`timescale 1ps/1ps
(* whitebox *)
module VCC (
    output wire VCC
);

    assign VCC = 1'b1;

endmodule
