module MULT25X18
  (
   A, B,
   OUT
   );

   input wire [24:0] A;
   input wire [17:0] B;

   output wire [85:0] OUT;

endmodule // MULT25X18

