(* blackbox *)
module LUT4 (I, O);
	input wire [3:0] I;
	output wire O;
endmodule
