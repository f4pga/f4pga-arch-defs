(* blackbox *)
module MULT (
	input [31:0] Amult,
	input [31:0] Bmult,
	input [1:0] Valid_mult,
	output [63:0] Cmult,
	input sel_mul_32x32
);

endmodule
