(* blackbox *)
module ASSP (
  input         WB_CLK,
  input         WBs_ACK,
  input  [31:0] WBs_RD_DAT,
  output [3:0]  WBs_BYTE_STB,
  output        WBs_CYC,
  output        WBs_WE,
  output        WBs_RD,
  output        WBs_STB,
  output [16:0] WBs_ADR,
  input  [3:0]  SDMA_Req,
  input  [3:0]  SDMA_Sreq,
  output [3:0]  SDMA_Done,
  output [3:0]  SDMA_Active,
  input  [3:0]  FB_msg_out,
  input  [7:0]  FB_Int_Clr,
  output        FB_Start,
  input         FB_Busy,
  output        WB_RST,
  output        Sys_PKfb_Rst,
  output        Sys_Clk0,
  output        Sys_Clk0_Rst,
  output        Sys_Clk1,
  output        Sys_Clk1_Rst,
  output        Sys_Pclk,
  output        Sys_Pclk_Rst,
  input         Sys_PKfb_Clk,
  input  [31:0] FB_PKfbData,
  output [31:0] WBs_WR_DAT,
  input  [3:0]  FB_PKfbPush,
  input         FB_PKfbSOF,
  input         FB_PKfbEOF,
  output [7:0]  Sensor_Int,
  output        FB_PKfbOverflow,
  output [23:0] TimeStamp,
  input         Sys_PSel,
  input  [15:0] SPIm_Paddr,
  input         SPIm_PEnable,
  input         SPIm_PWrite,
  input  [31:0] SPIm_PWdata,
  output        SPIm_PReady,
  output        SPIm_PSlvErr,
  output [31:0] SPIm_Prdata,
  input  [15:0] Device_ID,
  input  [13:0] FBIO_In_En,
  input  [13:0] FBIO_Out,
  input  [13:0] FBIO_Out_En,
  output [13:0] FBIO_In,
  //inout  [13:0] SFBIO, // FIXME: These should be "inout" but cannot model it this way
  input         Device_ID_6S, 
  input         Device_ID_4S, 
  input         SPIm_PWdata_26S, 
  input         SPIm_PWdata_24S,  
  input         SPIm_PWdata_14S, 
  input         SPIm_PWdata_11S, 
  input         SPIm_PWdata_0S, 
  input         SPIm_Paddr_8S, 
  input         SPIm_Paddr_6S, 
  input         FB_PKfbPush_1S, 
  input         FB_PKfbData_31S, 
  input         FB_PKfbData_21S,
  input         FB_PKfbData_19S,
  input         FB_PKfbData_9S,
  input         FB_PKfbData_6S,
  input         Sys_PKfb_ClkS,
  input         FB_BusyS,
  input         WB_CLKS
);

endmodule
