`default_nettype none
module INV(input A, output Z);
	assign Z = !A;
endmodule
