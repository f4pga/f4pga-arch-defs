module top (
	input  btn,
	output LED3,
);
	assign LED3 = btn;
endmodule
