`timescale 1ns/10ps
(* whitebox *)
module MULT (
			Amult,
			Bmult,
			Valid_mult,
			Cmult,
			sel_mul_32x32
			);

	input wire  [31:0] Amult;
	input wire  [31:0] Bmult;
	input wire   [1:0] Valid_mult;
	(* DELAY_MATRIX_Amult="{iopath_Amult0_Cmult0} {iopath_Amult0_Cmult1} {iopath_Amult0_Cmult2} {iopath_Amult0_Cmult3} {iopath_Amult0_Cmult4} {iopath_Amult0_Cmult5} {iopath_Amult0_Cmult6} {iopath_Amult0_Cmult7} {iopath_Amult0_Cmult8} {iopath_Amult0_Cmult9} {iopath_Amult0_Cmult10} {iopath_Amult0_Cmult11} {iopath_Amult0_Cmult12} {iopath_Amult0_Cmult13} {iopath_Amult0_Cmult14} {iopath_Amult0_Cmult15} {iopath_Amult0_Cmult16} {iopath_Amult0_Cmult17} {iopath_Amult0_Cmult18} {iopath_Amult0_Cmult19} {iopath_Amult0_Cmult20} {iopath_Amult0_Cmult21} {iopath_Amult0_Cmult22} {iopath_Amult0_Cmult23} {iopath_Amult0_Cmult24} {iopath_Amult0_Cmult25} {iopath_Amult0_Cmult26} {iopath_Amult0_Cmult27} {iopath_Amult0_Cmult28} {iopath_Amult0_Cmult29} {iopath_Amult0_Cmult30} {iopath_Amult0_Cmult31} {iopath_Amult0_Cmult32} {iopath_Amult0_Cmult33} {iopath_Amult0_Cmult34} {iopath_Amult0_Cmult35} {iopath_Amult0_Cmult36} {iopath_Amult0_Cmult37} {iopath_Amult0_Cmult38} {iopath_Amult0_Cmult39} {iopath_Amult0_Cmult40} {iopath_Amult0_Cmult41} {iopath_Amult0_Cmult42} {iopath_Amult0_Cmult43} {iopath_Amult0_Cmult44} {iopath_Amult0_Cmult45} {iopath_Amult0_Cmult46} {iopath_Amult0_Cmult47} {iopath_Amult0_Cmult48} {iopath_Amult0_Cmult49} {iopath_Amult0_Cmult50} {iopath_Amult0_Cmult51} {iopath_Amult0_Cmult52} {iopath_Amult0_Cmult53} {iopath_Amult0_Cmult54} {iopath_Amult0_Cmult55} {iopath_Amult0_Cmult56} {iopath_Amult0_Cmult57} {iopath_Amult0_Cmult58} {iopath_Amult0_Cmult59} {iopath_Amult0_Cmult60} {iopath_Amult0_Cmult61} {iopath_Amult0_Cmult62} {iopath_Amult0_Cmult63} 0 {iopath_Amult1_Cmult1} {iopath_Amult1_Cmult2} {iopath_Amult1_Cmult3} {iopath_Amult1_Cmult4} {iopath_Amult1_Cmult5} {iopath_Amult1_Cmult6} {iopath_Amult1_Cmult7} {iopath_Amult1_Cmult8} {iopath_Amult1_Cmult9} {iopath_Amult1_Cmult10} {iopath_Amult1_Cmult11} {iopath_Amult1_Cmult12} {iopath_Amult1_Cmult13} {iopath_Amult1_Cmult14} {iopath_Amult1_Cmult15} {iopath_Amult1_Cmult16} {iopath_Amult1_Cmult17} {iopath_Amult1_Cmult18} {iopath_Amult1_Cmult19} {iopath_Amult1_Cmult20} {iopath_Amult1_Cmult21} {iopath_Amult1_Cmult22} {iopath_Amult1_Cmult23} {iopath_Amult1_Cmult24} {iopath_Amult1_Cmult25} {iopath_Amult1_Cmult26} {iopath_Amult1_Cmult27} {iopath_Amult1_Cmult28} {iopath_Amult1_Cmult29} {iopath_Amult1_Cmult30} {iopath_Amult1_Cmult31} {iopath_Amult1_Cmult32} {iopath_Amult1_Cmult33} {iopath_Amult1_Cmult34} {iopath_Amult1_Cmult35} {iopath_Amult1_Cmult36} {iopath_Amult1_Cmult37} {iopath_Amult1_Cmult38} {iopath_Amult1_Cmult39} {iopath_Amult1_Cmult40} {iopath_Amult1_Cmult41} {iopath_Amult1_Cmult42} {iopath_Amult1_Cmult43} {iopath_Amult1_Cmult44} {iopath_Amult1_Cmult45} {iopath_Amult1_Cmult46} {iopath_Amult1_Cmult47} {iopath_Amult1_Cmult48} {iopath_Amult1_Cmult49} {iopath_Amult1_Cmult50} {iopath_Amult1_Cmult51} {iopath_Amult1_Cmult52} {iopath_Amult1_Cmult53} {iopath_Amult1_Cmult54} {iopath_Amult1_Cmult55} {iopath_Amult1_Cmult56} {iopath_Amult1_Cmult57} {iopath_Amult1_Cmult58} {iopath_Amult1_Cmult59} {iopath_Amult1_Cmult60} {iopath_Amult1_Cmult61} {iopath_Amult1_Cmult62} {iopath_Amult1_Cmult63} 0 0 {iopath_Amult2_Cmult2} {iopath_Amult2_Cmult3} {iopath_Amult2_Cmult4} {iopath_Amult2_Cmult5} {iopath_Amult2_Cmult6} {iopath_Amult2_Cmult7} {iopath_Amult2_Cmult8} {iopath_Amult2_Cmult9} {iopath_Amult2_Cmult10} {iopath_Amult2_Cmult11} {iopath_Amult2_Cmult12} {iopath_Amult2_Cmult13} {iopath_Amult2_Cmult14} {iopath_Amult2_Cmult15} {iopath_Amult2_Cmult16} {iopath_Amult2_Cmult17} {iopath_Amult2_Cmult18} {iopath_Amult2_Cmult19} {iopath_Amult2_Cmult20} {iopath_Amult2_Cmult21} {iopath_Amult2_Cmult22} {iopath_Amult2_Cmult23} {iopath_Amult2_Cmult24} {iopath_Amult2_Cmult25} {iopath_Amult2_Cmult26} {iopath_Amult2_Cmult27} {iopath_Amult2_Cmult28} {iopath_Amult2_Cmult29} {iopath_Amult2_Cmult30} {iopath_Amult2_Cmult31} {iopath_Amult2_Cmult32} {iopath_Amult2_Cmult33} {iopath_Amult2_Cmult34} {iopath_Amult2_Cmult35} {iopath_Amult2_Cmult36} {iopath_Amult2_Cmult37} {iopath_Amult2_Cmult38} {iopath_Amult2_Cmult39} {iopath_Amult2_Cmult40} {iopath_Amult2_Cmult41} {iopath_Amult2_Cmult42} {iopath_Amult2_Cmult43} {iopath_Amult2_Cmult44} {iopath_Amult2_Cmult45} {iopath_Amult2_Cmult46} {iopath_Amult2_Cmult47} {iopath_Amult2_Cmult48} {iopath_Amult2_Cmult49} {iopath_Amult2_Cmult50} {iopath_Amult2_Cmult51} {iopath_Amult2_Cmult52} {iopath_Amult2_Cmult53} {iopath_Amult2_Cmult54} {iopath_Amult2_Cmult55} {iopath_Amult2_Cmult56} {iopath_Amult2_Cmult57} {iopath_Amult2_Cmult58} {iopath_Amult2_Cmult59} {iopath_Amult2_Cmult60} {iopath_Amult2_Cmult61} {iopath_Amult2_Cmult62} {iopath_Amult2_Cmult63} 0 0 0 {iopath_Amult3_Cmult3} {iopath_Amult3_Cmult4} {iopath_Amult3_Cmult5} {iopath_Amult3_Cmult6} {iopath_Amult3_Cmult7} {iopath_Amult3_Cmult8} {iopath_Amult3_Cmult9} {iopath_Amult3_Cmult10} {iopath_Amult3_Cmult11} {iopath_Amult3_Cmult12} {iopath_Amult3_Cmult13} {iopath_Amult3_Cmult14} {iopath_Amult3_Cmult15} {iopath_Amult3_Cmult16} {iopath_Amult3_Cmult17} {iopath_Amult3_Cmult18} {iopath_Amult3_Cmult19} {iopath_Amult3_Cmult20} {iopath_Amult3_Cmult21} {iopath_Amult3_Cmult22} {iopath_Amult3_Cmult23} {iopath_Amult3_Cmult24} {iopath_Amult3_Cmult25} {iopath_Amult3_Cmult26} {iopath_Amult3_Cmult27} {iopath_Amult3_Cmult28} {iopath_Amult3_Cmult29} {iopath_Amult3_Cmult30} {iopath_Amult3_Cmult31} {iopath_Amult3_Cmult32} {iopath_Amult3_Cmult33} {iopath_Amult3_Cmult34} {iopath_Amult3_Cmult35} {iopath_Amult3_Cmult36} {iopath_Amult3_Cmult37} {iopath_Amult3_Cmult38} {iopath_Amult3_Cmult39} {iopath_Amult3_Cmult40} {iopath_Amult3_Cmult41} {iopath_Amult3_Cmult42} {iopath_Amult3_Cmult43} {iopath_Amult3_Cmult44} {iopath_Amult3_Cmult45} {iopath_Amult3_Cmult46} {iopath_Amult3_Cmult47} {iopath_Amult3_Cmult48} {iopath_Amult3_Cmult49} {iopath_Amult3_Cmult50} {iopath_Amult3_Cmult51} {iopath_Amult3_Cmult52} {iopath_Amult3_Cmult53} {iopath_Amult3_Cmult54} {iopath_Amult3_Cmult55} {iopath_Amult3_Cmult56} {iopath_Amult3_Cmult57} {iopath_Amult3_Cmult58} {iopath_Amult3_Cmult59} {iopath_Amult3_Cmult60} {iopath_Amult3_Cmult61} {iopath_Amult3_Cmult62} {iopath_Amult3_Cmult63} 0 0 0 0 {iopath_Amult4_Cmult4} {iopath_Amult4_Cmult5} {iopath_Amult4_Cmult6} {iopath_Amult4_Cmult7} {iopath_Amult4_Cmult8} {iopath_Amult4_Cmult9} {iopath_Amult4_Cmult10} {iopath_Amult4_Cmult11} {iopath_Amult4_Cmult12} {iopath_Amult4_Cmult13} {iopath_Amult4_Cmult14} {iopath_Amult4_Cmult15} {iopath_Amult4_Cmult16} {iopath_Amult4_Cmult17} {iopath_Amult4_Cmult18} {iopath_Amult4_Cmult19} {iopath_Amult4_Cmult20} {iopath_Amult4_Cmult21} {iopath_Amult4_Cmult22} {iopath_Amult4_Cmult23} {iopath_Amult4_Cmult24} {iopath_Amult4_Cmult25} {iopath_Amult4_Cmult26} {iopath_Amult4_Cmult27} {iopath_Amult4_Cmult28} {iopath_Amult4_Cmult29} {iopath_Amult4_Cmult30} {iopath_Amult4_Cmult31} {iopath_Amult4_Cmult32} {iopath_Amult4_Cmult33} {iopath_Amult4_Cmult34} {iopath_Amult4_Cmult35} {iopath_Amult4_Cmult36} {iopath_Amult4_Cmult37} {iopath_Amult4_Cmult38} {iopath_Amult4_Cmult39} {iopath_Amult4_Cmult40} {iopath_Amult4_Cmult41} {iopath_Amult4_Cmult42} {iopath_Amult4_Cmult43} {iopath_Amult4_Cmult44} {iopath_Amult4_Cmult45} {iopath_Amult4_Cmult46} {iopath_Amult4_Cmult47} {iopath_Amult4_Cmult48} {iopath_Amult4_Cmult49} {iopath_Amult4_Cmult50} {iopath_Amult4_Cmult51} {iopath_Amult4_Cmult52} {iopath_Amult4_Cmult53} {iopath_Amult4_Cmult54} {iopath_Amult4_Cmult55} {iopath_Amult4_Cmult56} {iopath_Amult4_Cmult57} {iopath_Amult4_Cmult58} {iopath_Amult4_Cmult59} {iopath_Amult4_Cmult60} {iopath_Amult4_Cmult61} {iopath_Amult4_Cmult62} {iopath_Amult4_Cmult63} 0 0 0 0 0 {iopath_Amult5_Cmult5} {iopath_Amult5_Cmult6} {iopath_Amult5_Cmult7} {iopath_Amult5_Cmult8} {iopath_Amult5_Cmult9} {iopath_Amult5_Cmult10} {iopath_Amult5_Cmult11} {iopath_Amult5_Cmult12} {iopath_Amult5_Cmult13} {iopath_Amult5_Cmult14} {iopath_Amult5_Cmult15} {iopath_Amult5_Cmult16} {iopath_Amult5_Cmult17} {iopath_Amult5_Cmult18} {iopath_Amult5_Cmult19} {iopath_Amult5_Cmult20} {iopath_Amult5_Cmult21} {iopath_Amult5_Cmult22} {iopath_Amult5_Cmult23} {iopath_Amult5_Cmult24} {iopath_Amult5_Cmult25} {iopath_Amult5_Cmult26} {iopath_Amult5_Cmult27} {iopath_Amult5_Cmult28} {iopath_Amult5_Cmult29} {iopath_Amult5_Cmult30} {iopath_Amult5_Cmult31} {iopath_Amult5_Cmult32} {iopath_Amult5_Cmult33} {iopath_Amult5_Cmult34} {iopath_Amult5_Cmult35} {iopath_Amult5_Cmult36} {iopath_Amult5_Cmult37} {iopath_Amult5_Cmult38} {iopath_Amult5_Cmult39} {iopath_Amult5_Cmult40} {iopath_Amult5_Cmult41} {iopath_Amult5_Cmult42} {iopath_Amult5_Cmult43} {iopath_Amult5_Cmult44} {iopath_Amult5_Cmult45} {iopath_Amult5_Cmult46} {iopath_Amult5_Cmult47} {iopath_Amult5_Cmult48} {iopath_Amult5_Cmult49} {iopath_Amult5_Cmult50} {iopath_Amult5_Cmult51} {iopath_Amult5_Cmult52} {iopath_Amult5_Cmult53} {iopath_Amult5_Cmult54} {iopath_Amult5_Cmult55} {iopath_Amult5_Cmult56} {iopath_Amult5_Cmult57} {iopath_Amult5_Cmult58} {iopath_Amult5_Cmult59} {iopath_Amult5_Cmult60} {iopath_Amult5_Cmult61} {iopath_Amult5_Cmult62} {iopath_Amult5_Cmult63} 0 0 0 0 0 0 {iopath_Amult6_Cmult6} {iopath_Amult6_Cmult7} {iopath_Amult6_Cmult8} {iopath_Amult6_Cmult9} {iopath_Amult6_Cmult10} {iopath_Amult6_Cmult11} {iopath_Amult6_Cmult12} {iopath_Amult6_Cmult13} {iopath_Amult6_Cmult14} {iopath_Amult6_Cmult15} {iopath_Amult6_Cmult16} {iopath_Amult6_Cmult17} {iopath_Amult6_Cmult18} {iopath_Amult6_Cmult19} {iopath_Amult6_Cmult20} {iopath_Amult6_Cmult21} {iopath_Amult6_Cmult22} {iopath_Amult6_Cmult23} {iopath_Amult6_Cmult24} {iopath_Amult6_Cmult25} {iopath_Amult6_Cmult26} {iopath_Amult6_Cmult27} {iopath_Amult6_Cmult28} {iopath_Amult6_Cmult29} {iopath_Amult6_Cmult30} {iopath_Amult6_Cmult31} {iopath_Amult6_Cmult32} {iopath_Amult6_Cmult33} {iopath_Amult6_Cmult34} {iopath_Amult6_Cmult35} {iopath_Amult6_Cmult36} {iopath_Amult6_Cmult37} {iopath_Amult6_Cmult38} {iopath_Amult6_Cmult39} {iopath_Amult6_Cmult40} {iopath_Amult6_Cmult41} {iopath_Amult6_Cmult42} {iopath_Amult6_Cmult43} {iopath_Amult6_Cmult44} {iopath_Amult6_Cmult45} {iopath_Amult6_Cmult46} {iopath_Amult6_Cmult47} {iopath_Amult6_Cmult48} {iopath_Amult6_Cmult49} {iopath_Amult6_Cmult50} {iopath_Amult6_Cmult51} {iopath_Amult6_Cmult52} {iopath_Amult6_Cmult53} {iopath_Amult6_Cmult54} {iopath_Amult6_Cmult55} {iopath_Amult6_Cmult56} {iopath_Amult6_Cmult57} {iopath_Amult6_Cmult58} {iopath_Amult6_Cmult59} {iopath_Amult6_Cmult60} {iopath_Amult6_Cmult61} {iopath_Amult6_Cmult62} {iopath_Amult6_Cmult63} 0 0 0 0 0 0 0 {iopath_Amult7_Cmult7} {iopath_Amult7_Cmult8} {iopath_Amult7_Cmult9} {iopath_Amult7_Cmult10} {iopath_Amult7_Cmult11} {iopath_Amult7_Cmult12} {iopath_Amult7_Cmult13} {iopath_Amult7_Cmult14} {iopath_Amult7_Cmult15} {iopath_Amult7_Cmult16} {iopath_Amult7_Cmult17} {iopath_Amult7_Cmult18} {iopath_Amult7_Cmult19} {iopath_Amult7_Cmult20} {iopath_Amult7_Cmult21} {iopath_Amult7_Cmult22} {iopath_Amult7_Cmult23} {iopath_Amult7_Cmult24} {iopath_Amult7_Cmult25} {iopath_Amult7_Cmult26} {iopath_Amult7_Cmult27} {iopath_Amult7_Cmult28} {iopath_Amult7_Cmult29} {iopath_Amult7_Cmult30} {iopath_Amult7_Cmult31} {iopath_Amult7_Cmult32} {iopath_Amult7_Cmult33} {iopath_Amult7_Cmult34} {iopath_Amult7_Cmult35} {iopath_Amult7_Cmult36} {iopath_Amult7_Cmult37} {iopath_Amult7_Cmult38} {iopath_Amult7_Cmult39} {iopath_Amult7_Cmult40} {iopath_Amult7_Cmult41} {iopath_Amult7_Cmult42} {iopath_Amult7_Cmult43} {iopath_Amult7_Cmult44} {iopath_Amult7_Cmult45} {iopath_Amult7_Cmult46} {iopath_Amult7_Cmult47} {iopath_Amult7_Cmult48} {iopath_Amult7_Cmult49} {iopath_Amult7_Cmult50} {iopath_Amult7_Cmult51} {iopath_Amult7_Cmult52} {iopath_Amult7_Cmult53} {iopath_Amult7_Cmult54} {iopath_Amult7_Cmult55} {iopath_Amult7_Cmult56} {iopath_Amult7_Cmult57} {iopath_Amult7_Cmult58} {iopath_Amult7_Cmult59} {iopath_Amult7_Cmult60} {iopath_Amult7_Cmult61} {iopath_Amult7_Cmult62} {iopath_Amult7_Cmult63} 0 0 0 0 0 0 0 0 {iopath_Amult8_Cmult8} {iopath_Amult8_Cmult9} {iopath_Amult8_Cmult10} {iopath_Amult8_Cmult11} {iopath_Amult8_Cmult12} {iopath_Amult8_Cmult13} {iopath_Amult8_Cmult14} {iopath_Amult8_Cmult15} {iopath_Amult8_Cmult16} {iopath_Amult8_Cmult17} {iopath_Amult8_Cmult18} {iopath_Amult8_Cmult19} {iopath_Amult8_Cmult20} {iopath_Amult8_Cmult21} {iopath_Amult8_Cmult22} {iopath_Amult8_Cmult23} {iopath_Amult8_Cmult24} {iopath_Amult8_Cmult25} {iopath_Amult8_Cmult26} {iopath_Amult8_Cmult27} {iopath_Amult8_Cmult28} {iopath_Amult8_Cmult29} {iopath_Amult8_Cmult30} {iopath_Amult8_Cmult31} {iopath_Amult8_Cmult32} {iopath_Amult8_Cmult33} {iopath_Amult8_Cmult34} {iopath_Amult8_Cmult35} {iopath_Amult8_Cmult36} {iopath_Amult8_Cmult37} {iopath_Amult8_Cmult38} {iopath_Amult8_Cmult39} {iopath_Amult8_Cmult40} {iopath_Amult8_Cmult41} {iopath_Amult8_Cmult42} {iopath_Amult8_Cmult43} {iopath_Amult8_Cmult44} {iopath_Amult8_Cmult45} {iopath_Amult8_Cmult46} {iopath_Amult8_Cmult47} {iopath_Amult8_Cmult48} {iopath_Amult8_Cmult49} {iopath_Amult8_Cmult50} {iopath_Amult8_Cmult51} {iopath_Amult8_Cmult52} {iopath_Amult8_Cmult53} {iopath_Amult8_Cmult54} {iopath_Amult8_Cmult55} {iopath_Amult8_Cmult56} {iopath_Amult8_Cmult57} {iopath_Amult8_Cmult58} {iopath_Amult8_Cmult59} {iopath_Amult8_Cmult60} {iopath_Amult8_Cmult61} {iopath_Amult8_Cmult62} {iopath_Amult8_Cmult63} 0 0 0 0 0 0 0 0 0 {iopath_Amult9_Cmult9} {iopath_Amult9_Cmult10} {iopath_Amult9_Cmult11} {iopath_Amult9_Cmult12} {iopath_Amult9_Cmult13} {iopath_Amult9_Cmult14} {iopath_Amult9_Cmult15} {iopath_Amult9_Cmult16} {iopath_Amult9_Cmult17} {iopath_Amult9_Cmult18} {iopath_Amult9_Cmult19} {iopath_Amult9_Cmult20} {iopath_Amult9_Cmult21} {iopath_Amult9_Cmult22} {iopath_Amult9_Cmult23} {iopath_Amult9_Cmult24} {iopath_Amult9_Cmult25} {iopath_Amult9_Cmult26} {iopath_Amult9_Cmult27} {iopath_Amult9_Cmult28} {iopath_Amult9_Cmult29} {iopath_Amult9_Cmult30} {iopath_Amult9_Cmult31} {iopath_Amult9_Cmult32} {iopath_Amult9_Cmult33} {iopath_Amult9_Cmult34} {iopath_Amult9_Cmult35} {iopath_Amult9_Cmult36} {iopath_Amult9_Cmult37} {iopath_Amult9_Cmult38} {iopath_Amult9_Cmult39} {iopath_Amult9_Cmult40} {iopath_Amult9_Cmult41} {iopath_Amult9_Cmult42} {iopath_Amult9_Cmult43} {iopath_Amult9_Cmult44} {iopath_Amult9_Cmult45} {iopath_Amult9_Cmult46} {iopath_Amult9_Cmult47} {iopath_Amult9_Cmult48} {iopath_Amult9_Cmult49} {iopath_Amult9_Cmult50} {iopath_Amult9_Cmult51} {iopath_Amult9_Cmult52} {iopath_Amult9_Cmult53} {iopath_Amult9_Cmult54} {iopath_Amult9_Cmult55} {iopath_Amult9_Cmult56} {iopath_Amult9_Cmult57} {iopath_Amult9_Cmult58} {iopath_Amult9_Cmult59} {iopath_Amult9_Cmult60} {iopath_Amult9_Cmult61} {iopath_Amult9_Cmult62} {iopath_Amult9_Cmult63} 0 0 0 0 0 0 0 0 0 0 {iopath_Amult10_Cmult10} {iopath_Amult10_Cmult11} {iopath_Amult10_Cmult12} {iopath_Amult10_Cmult13} {iopath_Amult10_Cmult14} {iopath_Amult10_Cmult15} {iopath_Amult10_Cmult16} {iopath_Amult10_Cmult17} {iopath_Amult10_Cmult18} {iopath_Amult10_Cmult19} {iopath_Amult10_Cmult20} {iopath_Amult10_Cmult21} {iopath_Amult10_Cmult22} {iopath_Amult10_Cmult23} {iopath_Amult10_Cmult24} {iopath_Amult10_Cmult25} {iopath_Amult10_Cmult26} {iopath_Amult10_Cmult27} {iopath_Amult10_Cmult28} {iopath_Amult10_Cmult29} {iopath_Amult10_Cmult30} {iopath_Amult10_Cmult31} {iopath_Amult10_Cmult32} {iopath_Amult10_Cmult33} {iopath_Amult10_Cmult34} {iopath_Amult10_Cmult35} {iopath_Amult10_Cmult36} {iopath_Amult10_Cmult37} {iopath_Amult10_Cmult38} {iopath_Amult10_Cmult39} {iopath_Amult10_Cmult40} {iopath_Amult10_Cmult41} {iopath_Amult10_Cmult42} {iopath_Amult10_Cmult43} {iopath_Amult10_Cmult44} {iopath_Amult10_Cmult45} {iopath_Amult10_Cmult46} {iopath_Amult10_Cmult47} {iopath_Amult10_Cmult48} {iopath_Amult10_Cmult49} {iopath_Amult10_Cmult50} {iopath_Amult10_Cmult51} {iopath_Amult10_Cmult52} {iopath_Amult10_Cmult53} {iopath_Amult10_Cmult54} {iopath_Amult10_Cmult55} {iopath_Amult10_Cmult56} {iopath_Amult10_Cmult57} {iopath_Amult10_Cmult58} {iopath_Amult10_Cmult59} {iopath_Amult10_Cmult60} {iopath_Amult10_Cmult61} {iopath_Amult10_Cmult62} {iopath_Amult10_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult11_Cmult11} {iopath_Amult11_Cmult12} {iopath_Amult11_Cmult13} {iopath_Amult11_Cmult14} {iopath_Amult11_Cmult15} {iopath_Amult11_Cmult16} {iopath_Amult11_Cmult17} {iopath_Amult11_Cmult18} {iopath_Amult11_Cmult19} {iopath_Amult11_Cmult20} {iopath_Amult11_Cmult21} {iopath_Amult11_Cmult22} {iopath_Amult11_Cmult23} {iopath_Amult11_Cmult24} {iopath_Amult11_Cmult25} {iopath_Amult11_Cmult26} {iopath_Amult11_Cmult27} {iopath_Amult11_Cmult28} {iopath_Amult11_Cmult29} {iopath_Amult11_Cmult30} {iopath_Amult11_Cmult31} {iopath_Amult11_Cmult32} {iopath_Amult11_Cmult33} {iopath_Amult11_Cmult34} {iopath_Amult11_Cmult35} {iopath_Amult11_Cmult36} {iopath_Amult11_Cmult37} {iopath_Amult11_Cmult38} {iopath_Amult11_Cmult39} {iopath_Amult11_Cmult40} {iopath_Amult11_Cmult41} {iopath_Amult11_Cmult42} {iopath_Amult11_Cmult43} {iopath_Amult11_Cmult44} {iopath_Amult11_Cmult45} {iopath_Amult11_Cmult46} {iopath_Amult11_Cmult47} {iopath_Amult11_Cmult48} {iopath_Amult11_Cmult49} {iopath_Amult11_Cmult50} {iopath_Amult11_Cmult51} {iopath_Amult11_Cmult52} {iopath_Amult11_Cmult53} {iopath_Amult11_Cmult54} {iopath_Amult11_Cmult55} {iopath_Amult11_Cmult56} {iopath_Amult11_Cmult57} {iopath_Amult11_Cmult58} {iopath_Amult11_Cmult59} {iopath_Amult11_Cmult60} {iopath_Amult11_Cmult61} {iopath_Amult11_Cmult62} {iopath_Amult11_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult12_Cmult12} {iopath_Amult12_Cmult13} {iopath_Amult12_Cmult14} {iopath_Amult12_Cmult15} {iopath_Amult12_Cmult16} {iopath_Amult12_Cmult17} {iopath_Amult12_Cmult18} {iopath_Amult12_Cmult19} {iopath_Amult12_Cmult20} {iopath_Amult12_Cmult21} {iopath_Amult12_Cmult22} {iopath_Amult12_Cmult23} {iopath_Amult12_Cmult24} {iopath_Amult12_Cmult25} {iopath_Amult12_Cmult26} {iopath_Amult12_Cmult27} {iopath_Amult12_Cmult28} {iopath_Amult12_Cmult29} {iopath_Amult12_Cmult30} {iopath_Amult12_Cmult31} {iopath_Amult12_Cmult32} {iopath_Amult12_Cmult33} {iopath_Amult12_Cmult34} {iopath_Amult12_Cmult35} {iopath_Amult12_Cmult36} {iopath_Amult12_Cmult37} {iopath_Amult12_Cmult38} {iopath_Amult12_Cmult39} {iopath_Amult12_Cmult40} {iopath_Amult12_Cmult41} {iopath_Amult12_Cmult42} {iopath_Amult12_Cmult43} {iopath_Amult12_Cmult44} {iopath_Amult12_Cmult45} {iopath_Amult12_Cmult46} {iopath_Amult12_Cmult47} {iopath_Amult12_Cmult48} {iopath_Amult12_Cmult49} {iopath_Amult12_Cmult50} {iopath_Amult12_Cmult51} {iopath_Amult12_Cmult52} {iopath_Amult12_Cmult53} {iopath_Amult12_Cmult54} {iopath_Amult12_Cmult55} {iopath_Amult12_Cmult56} {iopath_Amult12_Cmult57} {iopath_Amult12_Cmult58} {iopath_Amult12_Cmult59} {iopath_Amult12_Cmult60} {iopath_Amult12_Cmult61} {iopath_Amult12_Cmult62} {iopath_Amult12_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult13_Cmult13} {iopath_Amult13_Cmult14} {iopath_Amult13_Cmult15} {iopath_Amult13_Cmult16} {iopath_Amult13_Cmult17} {iopath_Amult13_Cmult18} {iopath_Amult13_Cmult19} {iopath_Amult13_Cmult20} {iopath_Amult13_Cmult21} {iopath_Amult13_Cmult22} {iopath_Amult13_Cmult23} {iopath_Amult13_Cmult24} {iopath_Amult13_Cmult25} {iopath_Amult13_Cmult26} {iopath_Amult13_Cmult27} {iopath_Amult13_Cmult28} {iopath_Amult13_Cmult29} {iopath_Amult13_Cmult30} {iopath_Amult13_Cmult31} {iopath_Amult13_Cmult32} {iopath_Amult13_Cmult33} {iopath_Amult13_Cmult34} {iopath_Amult13_Cmult35} {iopath_Amult13_Cmult36} {iopath_Amult13_Cmult37} {iopath_Amult13_Cmult38} {iopath_Amult13_Cmult39} {iopath_Amult13_Cmult40} {iopath_Amult13_Cmult41} {iopath_Amult13_Cmult42} {iopath_Amult13_Cmult43} {iopath_Amult13_Cmult44} {iopath_Amult13_Cmult45} {iopath_Amult13_Cmult46} {iopath_Amult13_Cmult47} {iopath_Amult13_Cmult48} {iopath_Amult13_Cmult49} {iopath_Amult13_Cmult50} {iopath_Amult13_Cmult51} {iopath_Amult13_Cmult52} {iopath_Amult13_Cmult53} {iopath_Amult13_Cmult54} {iopath_Amult13_Cmult55} {iopath_Amult13_Cmult56} {iopath_Amult13_Cmult57} {iopath_Amult13_Cmult58} {iopath_Amult13_Cmult59} {iopath_Amult13_Cmult60} {iopath_Amult13_Cmult61} {iopath_Amult13_Cmult62} {iopath_Amult13_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult14_Cmult14} {iopath_Amult14_Cmult15} {iopath_Amult14_Cmult16} {iopath_Amult14_Cmult17} {iopath_Amult14_Cmult18} {iopath_Amult14_Cmult19} {iopath_Amult14_Cmult20} {iopath_Amult14_Cmult21} {iopath_Amult14_Cmult22} {iopath_Amult14_Cmult23} {iopath_Amult14_Cmult24} {iopath_Amult14_Cmult25} {iopath_Amult14_Cmult26} {iopath_Amult14_Cmult27} {iopath_Amult14_Cmult28} {iopath_Amult14_Cmult29} {iopath_Amult14_Cmult30} {iopath_Amult14_Cmult31} {iopath_Amult14_Cmult32} {iopath_Amult14_Cmult33} {iopath_Amult14_Cmult34} {iopath_Amult14_Cmult35} {iopath_Amult14_Cmult36} {iopath_Amult14_Cmult37} {iopath_Amult14_Cmult38} {iopath_Amult14_Cmult39} {iopath_Amult14_Cmult40} {iopath_Amult14_Cmult41} {iopath_Amult14_Cmult42} {iopath_Amult14_Cmult43} {iopath_Amult14_Cmult44} {iopath_Amult14_Cmult45} {iopath_Amult14_Cmult46} {iopath_Amult14_Cmult47} {iopath_Amult14_Cmult48} {iopath_Amult14_Cmult49} {iopath_Amult14_Cmult50} {iopath_Amult14_Cmult51} {iopath_Amult14_Cmult52} {iopath_Amult14_Cmult53} {iopath_Amult14_Cmult54} {iopath_Amult14_Cmult55} {iopath_Amult14_Cmult56} {iopath_Amult14_Cmult57} {iopath_Amult14_Cmult58} {iopath_Amult14_Cmult59} {iopath_Amult14_Cmult60} {iopath_Amult14_Cmult61} {iopath_Amult14_Cmult62} {iopath_Amult14_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult15_Cmult15} {iopath_Amult15_Cmult16} {iopath_Amult15_Cmult17} {iopath_Amult15_Cmult18} {iopath_Amult15_Cmult19} {iopath_Amult15_Cmult20} {iopath_Amult15_Cmult21} {iopath_Amult15_Cmult22} {iopath_Amult15_Cmult23} {iopath_Amult15_Cmult24} {iopath_Amult15_Cmult25} {iopath_Amult15_Cmult26} {iopath_Amult15_Cmult27} {iopath_Amult15_Cmult28} {iopath_Amult15_Cmult29} {iopath_Amult15_Cmult30} {iopath_Amult15_Cmult31} {iopath_Amult15_Cmult32} {iopath_Amult15_Cmult33} {iopath_Amult15_Cmult34} {iopath_Amult15_Cmult35} {iopath_Amult15_Cmult36} {iopath_Amult15_Cmult37} {iopath_Amult15_Cmult38} {iopath_Amult15_Cmult39} {iopath_Amult15_Cmult40} {iopath_Amult15_Cmult41} {iopath_Amult15_Cmult42} {iopath_Amult15_Cmult43} {iopath_Amult15_Cmult44} {iopath_Amult15_Cmult45} {iopath_Amult15_Cmult46} {iopath_Amult15_Cmult47} {iopath_Amult15_Cmult48} {iopath_Amult15_Cmult49} {iopath_Amult15_Cmult50} {iopath_Amult15_Cmult51} {iopath_Amult15_Cmult52} {iopath_Amult15_Cmult53} {iopath_Amult15_Cmult54} {iopath_Amult15_Cmult55} {iopath_Amult15_Cmult56} {iopath_Amult15_Cmult57} {iopath_Amult15_Cmult58} {iopath_Amult15_Cmult59} {iopath_Amult15_Cmult60} {iopath_Amult15_Cmult61} {iopath_Amult15_Cmult62} {iopath_Amult15_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult16_Cmult16} {iopath_Amult16_Cmult17} {iopath_Amult16_Cmult18} {iopath_Amult16_Cmult19} {iopath_Amult16_Cmult20} {iopath_Amult16_Cmult21} {iopath_Amult16_Cmult22} {iopath_Amult16_Cmult23} {iopath_Amult16_Cmult24} {iopath_Amult16_Cmult25} {iopath_Amult16_Cmult26} {iopath_Amult16_Cmult27} {iopath_Amult16_Cmult28} {iopath_Amult16_Cmult29} {iopath_Amult16_Cmult30} {iopath_Amult16_Cmult31} {iopath_Amult16_Cmult32} {iopath_Amult16_Cmult33} {iopath_Amult16_Cmult34} {iopath_Amult16_Cmult35} {iopath_Amult16_Cmult36} {iopath_Amult16_Cmult37} {iopath_Amult16_Cmult38} {iopath_Amult16_Cmult39} {iopath_Amult16_Cmult40} {iopath_Amult16_Cmult41} {iopath_Amult16_Cmult42} {iopath_Amult16_Cmult43} {iopath_Amult16_Cmult44} {iopath_Amult16_Cmult45} {iopath_Amult16_Cmult46} {iopath_Amult16_Cmult47} {iopath_Amult16_Cmult48} {iopath_Amult16_Cmult49} {iopath_Amult16_Cmult50} {iopath_Amult16_Cmult51} {iopath_Amult16_Cmult52} {iopath_Amult16_Cmult53} {iopath_Amult16_Cmult54} {iopath_Amult16_Cmult55} {iopath_Amult16_Cmult56} {iopath_Amult16_Cmult57} {iopath_Amult16_Cmult58} {iopath_Amult16_Cmult59} {iopath_Amult16_Cmult60} {iopath_Amult16_Cmult61} {iopath_Amult16_Cmult62} {iopath_Amult16_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult17_Cmult17} {iopath_Amult17_Cmult18} {iopath_Amult17_Cmult19} {iopath_Amult17_Cmult20} {iopath_Amult17_Cmult21} {iopath_Amult17_Cmult22} {iopath_Amult17_Cmult23} {iopath_Amult17_Cmult24} {iopath_Amult17_Cmult25} {iopath_Amult17_Cmult26} {iopath_Amult17_Cmult27} {iopath_Amult17_Cmult28} {iopath_Amult17_Cmult29} {iopath_Amult17_Cmult30} {iopath_Amult17_Cmult31} {iopath_Amult17_Cmult32} {iopath_Amult17_Cmult33} {iopath_Amult17_Cmult34} {iopath_Amult17_Cmult35} {iopath_Amult17_Cmult36} {iopath_Amult17_Cmult37} {iopath_Amult17_Cmult38} {iopath_Amult17_Cmult39} {iopath_Amult17_Cmult40} {iopath_Amult17_Cmult41} {iopath_Amult17_Cmult42} {iopath_Amult17_Cmult43} {iopath_Amult17_Cmult44} {iopath_Amult17_Cmult45} {iopath_Amult17_Cmult46} {iopath_Amult17_Cmult47} {iopath_Amult17_Cmult48} {iopath_Amult17_Cmult49} {iopath_Amult17_Cmult50} {iopath_Amult17_Cmult51} {iopath_Amult17_Cmult52} {iopath_Amult17_Cmult53} {iopath_Amult17_Cmult54} {iopath_Amult17_Cmult55} {iopath_Amult17_Cmult56} {iopath_Amult17_Cmult57} {iopath_Amult17_Cmult58} {iopath_Amult17_Cmult59} {iopath_Amult17_Cmult60} {iopath_Amult17_Cmult61} {iopath_Amult17_Cmult62} {iopath_Amult17_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult18_Cmult18} {iopath_Amult18_Cmult19} {iopath_Amult18_Cmult20} {iopath_Amult18_Cmult21} {iopath_Amult18_Cmult22} {iopath_Amult18_Cmult23} {iopath_Amult18_Cmult24} {iopath_Amult18_Cmult25} {iopath_Amult18_Cmult26} {iopath_Amult18_Cmult27} {iopath_Amult18_Cmult28} {iopath_Amult18_Cmult29} {iopath_Amult18_Cmult30} {iopath_Amult18_Cmult31} {iopath_Amult18_Cmult32} {iopath_Amult18_Cmult33} {iopath_Amult18_Cmult34} {iopath_Amult18_Cmult35} {iopath_Amult18_Cmult36} {iopath_Amult18_Cmult37} {iopath_Amult18_Cmult38} {iopath_Amult18_Cmult39} {iopath_Amult18_Cmult40} {iopath_Amult18_Cmult41} {iopath_Amult18_Cmult42} {iopath_Amult18_Cmult43} {iopath_Amult18_Cmult44} {iopath_Amult18_Cmult45} {iopath_Amult18_Cmult46} {iopath_Amult18_Cmult47} {iopath_Amult18_Cmult48} {iopath_Amult18_Cmult49} {iopath_Amult18_Cmult50} {iopath_Amult18_Cmult51} {iopath_Amult18_Cmult52} {iopath_Amult18_Cmult53} {iopath_Amult18_Cmult54} {iopath_Amult18_Cmult55} {iopath_Amult18_Cmult56} {iopath_Amult18_Cmult57} {iopath_Amult18_Cmult58} {iopath_Amult18_Cmult59} {iopath_Amult18_Cmult60} {iopath_Amult18_Cmult61} {iopath_Amult18_Cmult62} {iopath_Amult18_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult19_Cmult19} {iopath_Amult19_Cmult20} {iopath_Amult19_Cmult21} {iopath_Amult19_Cmult22} {iopath_Amult19_Cmult23} {iopath_Amult19_Cmult24} {iopath_Amult19_Cmult25} {iopath_Amult19_Cmult26} {iopath_Amult19_Cmult27} {iopath_Amult19_Cmult28} {iopath_Amult19_Cmult29} {iopath_Amult19_Cmult30} {iopath_Amult19_Cmult31} {iopath_Amult19_Cmult32} {iopath_Amult19_Cmult33} {iopath_Amult19_Cmult34} {iopath_Amult19_Cmult35} {iopath_Amult19_Cmult36} {iopath_Amult19_Cmult37} {iopath_Amult19_Cmult38} {iopath_Amult19_Cmult39} {iopath_Amult19_Cmult40} {iopath_Amult19_Cmult41} {iopath_Amult19_Cmult42} {iopath_Amult19_Cmult43} {iopath_Amult19_Cmult44} {iopath_Amult19_Cmult45} {iopath_Amult19_Cmult46} {iopath_Amult19_Cmult47} {iopath_Amult19_Cmult48} {iopath_Amult19_Cmult49} {iopath_Amult19_Cmult50} {iopath_Amult19_Cmult51} {iopath_Amult19_Cmult52} {iopath_Amult19_Cmult53} {iopath_Amult19_Cmult54} {iopath_Amult19_Cmult55} {iopath_Amult19_Cmult56} {iopath_Amult19_Cmult57} {iopath_Amult19_Cmult58} {iopath_Amult19_Cmult59} {iopath_Amult19_Cmult60} {iopath_Amult19_Cmult61} {iopath_Amult19_Cmult62} {iopath_Amult19_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult20_Cmult20} {iopath_Amult20_Cmult21} {iopath_Amult20_Cmult22} {iopath_Amult20_Cmult23} {iopath_Amult20_Cmult24} {iopath_Amult20_Cmult25} {iopath_Amult20_Cmult26} {iopath_Amult20_Cmult27} {iopath_Amult20_Cmult28} {iopath_Amult20_Cmult29} {iopath_Amult20_Cmult30} {iopath_Amult20_Cmult31} {iopath_Amult20_Cmult32} {iopath_Amult20_Cmult33} {iopath_Amult20_Cmult34} {iopath_Amult20_Cmult35} {iopath_Amult20_Cmult36} {iopath_Amult20_Cmult37} {iopath_Amult20_Cmult38} {iopath_Amult20_Cmult39} {iopath_Amult20_Cmult40} {iopath_Amult20_Cmult41} {iopath_Amult20_Cmult42} {iopath_Amult20_Cmult43} {iopath_Amult20_Cmult44} {iopath_Amult20_Cmult45} {iopath_Amult20_Cmult46} {iopath_Amult20_Cmult47} {iopath_Amult20_Cmult48} {iopath_Amult20_Cmult49} {iopath_Amult20_Cmult50} {iopath_Amult20_Cmult51} {iopath_Amult20_Cmult52} {iopath_Amult20_Cmult53} {iopath_Amult20_Cmult54} {iopath_Amult20_Cmult55} {iopath_Amult20_Cmult56} {iopath_Amult20_Cmult57} {iopath_Amult20_Cmult58} {iopath_Amult20_Cmult59} {iopath_Amult20_Cmult60} {iopath_Amult20_Cmult61} {iopath_Amult20_Cmult62} {iopath_Amult20_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult21_Cmult21} {iopath_Amult21_Cmult22} {iopath_Amult21_Cmult23} {iopath_Amult21_Cmult24} {iopath_Amult21_Cmult25} {iopath_Amult21_Cmult26} {iopath_Amult21_Cmult27} {iopath_Amult21_Cmult28} {iopath_Amult21_Cmult29} {iopath_Amult21_Cmult30} {iopath_Amult21_Cmult31} {iopath_Amult21_Cmult32} {iopath_Amult21_Cmult33} {iopath_Amult21_Cmult34} {iopath_Amult21_Cmult35} {iopath_Amult21_Cmult36} {iopath_Amult21_Cmult37} {iopath_Amult21_Cmult38} {iopath_Amult21_Cmult39} {iopath_Amult21_Cmult40} {iopath_Amult21_Cmult41} {iopath_Amult21_Cmult42} {iopath_Amult21_Cmult43} {iopath_Amult21_Cmult44} {iopath_Amult21_Cmult45} {iopath_Amult21_Cmult46} {iopath_Amult21_Cmult47} {iopath_Amult21_Cmult48} {iopath_Amult21_Cmult49} {iopath_Amult21_Cmult50} {iopath_Amult21_Cmult51} {iopath_Amult21_Cmult52} {iopath_Amult21_Cmult53} {iopath_Amult21_Cmult54} {iopath_Amult21_Cmult55} {iopath_Amult21_Cmult56} {iopath_Amult21_Cmult57} {iopath_Amult21_Cmult58} {iopath_Amult21_Cmult59} {iopath_Amult21_Cmult60} {iopath_Amult21_Cmult61} {iopath_Amult21_Cmult62} {iopath_Amult21_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult22_Cmult22} {iopath_Amult22_Cmult23} {iopath_Amult22_Cmult24} {iopath_Amult22_Cmult25} {iopath_Amult22_Cmult26} {iopath_Amult22_Cmult27} {iopath_Amult22_Cmult28} {iopath_Amult22_Cmult29} {iopath_Amult22_Cmult30} {iopath_Amult22_Cmult31} {iopath_Amult22_Cmult32} {iopath_Amult22_Cmult33} {iopath_Amult22_Cmult34} {iopath_Amult22_Cmult35} {iopath_Amult22_Cmult36} {iopath_Amult22_Cmult37} {iopath_Amult22_Cmult38} {iopath_Amult22_Cmult39} {iopath_Amult22_Cmult40} {iopath_Amult22_Cmult41} {iopath_Amult22_Cmult42} {iopath_Amult22_Cmult43} {iopath_Amult22_Cmult44} {iopath_Amult22_Cmult45} {iopath_Amult22_Cmult46} {iopath_Amult22_Cmult47} {iopath_Amult22_Cmult48} {iopath_Amult22_Cmult49} {iopath_Amult22_Cmult50} {iopath_Amult22_Cmult51} {iopath_Amult22_Cmult52} {iopath_Amult22_Cmult53} {iopath_Amult22_Cmult54} {iopath_Amult22_Cmult55} {iopath_Amult22_Cmult56} {iopath_Amult22_Cmult57} {iopath_Amult22_Cmult58} {iopath_Amult22_Cmult59} {iopath_Amult22_Cmult60} {iopath_Amult22_Cmult61} {iopath_Amult22_Cmult62} {iopath_Amult22_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult23_Cmult23} {iopath_Amult23_Cmult24} {iopath_Amult23_Cmult25} {iopath_Amult23_Cmult26} {iopath_Amult23_Cmult27} {iopath_Amult23_Cmult28} {iopath_Amult23_Cmult29} {iopath_Amult23_Cmult30} {iopath_Amult23_Cmult31} {iopath_Amult23_Cmult32} {iopath_Amult23_Cmult33} {iopath_Amult23_Cmult34} {iopath_Amult23_Cmult35} {iopath_Amult23_Cmult36} {iopath_Amult23_Cmult37} {iopath_Amult23_Cmult38} {iopath_Amult23_Cmult39} {iopath_Amult23_Cmult40} {iopath_Amult23_Cmult41} {iopath_Amult23_Cmult42} {iopath_Amult23_Cmult43} {iopath_Amult23_Cmult44} {iopath_Amult23_Cmult45} {iopath_Amult23_Cmult46} {iopath_Amult23_Cmult47} {iopath_Amult23_Cmult48} {iopath_Amult23_Cmult49} {iopath_Amult23_Cmult50} {iopath_Amult23_Cmult51} {iopath_Amult23_Cmult52} {iopath_Amult23_Cmult53} {iopath_Amult23_Cmult54} {iopath_Amult23_Cmult55} {iopath_Amult23_Cmult56} {iopath_Amult23_Cmult57} {iopath_Amult23_Cmult58} {iopath_Amult23_Cmult59} {iopath_Amult23_Cmult60} {iopath_Amult23_Cmult61} {iopath_Amult23_Cmult62} {iopath_Amult23_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult24_Cmult24} {iopath_Amult24_Cmult25} {iopath_Amult24_Cmult26} {iopath_Amult24_Cmult27} {iopath_Amult24_Cmult28} {iopath_Amult24_Cmult29} {iopath_Amult24_Cmult30} {iopath_Amult24_Cmult31} {iopath_Amult24_Cmult32} {iopath_Amult24_Cmult33} {iopath_Amult24_Cmult34} {iopath_Amult24_Cmult35} {iopath_Amult24_Cmult36} {iopath_Amult24_Cmult37} {iopath_Amult24_Cmult38} {iopath_Amult24_Cmult39} {iopath_Amult24_Cmult40} {iopath_Amult24_Cmult41} {iopath_Amult24_Cmult42} {iopath_Amult24_Cmult43} {iopath_Amult24_Cmult44} {iopath_Amult24_Cmult45} {iopath_Amult24_Cmult46} {iopath_Amult24_Cmult47} {iopath_Amult24_Cmult48} {iopath_Amult24_Cmult49} {iopath_Amult24_Cmult50} {iopath_Amult24_Cmult51} {iopath_Amult24_Cmult52} {iopath_Amult24_Cmult53} {iopath_Amult24_Cmult54} {iopath_Amult24_Cmult55} {iopath_Amult24_Cmult56} {iopath_Amult24_Cmult57} {iopath_Amult24_Cmult58} {iopath_Amult24_Cmult59} {iopath_Amult24_Cmult60} {iopath_Amult24_Cmult61} {iopath_Amult24_Cmult62} {iopath_Amult24_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult25_Cmult25} {iopath_Amult25_Cmult26} {iopath_Amult25_Cmult27} {iopath_Amult25_Cmult28} {iopath_Amult25_Cmult29} {iopath_Amult25_Cmult30} {iopath_Amult25_Cmult31} {iopath_Amult25_Cmult32} {iopath_Amult25_Cmult33} {iopath_Amult25_Cmult34} {iopath_Amult25_Cmult35} {iopath_Amult25_Cmult36} {iopath_Amult25_Cmult37} {iopath_Amult25_Cmult38} {iopath_Amult25_Cmult39} {iopath_Amult25_Cmult40} {iopath_Amult25_Cmult41} {iopath_Amult25_Cmult42} {iopath_Amult25_Cmult43} {iopath_Amult25_Cmult44} {iopath_Amult25_Cmult45} {iopath_Amult25_Cmult46} {iopath_Amult25_Cmult47} {iopath_Amult25_Cmult48} {iopath_Amult25_Cmult49} {iopath_Amult25_Cmult50} {iopath_Amult25_Cmult51} {iopath_Amult25_Cmult52} {iopath_Amult25_Cmult53} {iopath_Amult25_Cmult54} {iopath_Amult25_Cmult55} {iopath_Amult25_Cmult56} {iopath_Amult25_Cmult57} {iopath_Amult25_Cmult58} {iopath_Amult25_Cmult59} {iopath_Amult25_Cmult60} {iopath_Amult25_Cmult61} {iopath_Amult25_Cmult62} {iopath_Amult25_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult26_Cmult26} {iopath_Amult26_Cmult27} {iopath_Amult26_Cmult28} {iopath_Amult26_Cmult29} {iopath_Amult26_Cmult30} {iopath_Amult26_Cmult31} {iopath_Amult26_Cmult32} {iopath_Amult26_Cmult33} {iopath_Amult26_Cmult34} {iopath_Amult26_Cmult35} {iopath_Amult26_Cmult36} {iopath_Amult26_Cmult37} {iopath_Amult26_Cmult38} {iopath_Amult26_Cmult39} {iopath_Amult26_Cmult40} {iopath_Amult26_Cmult41} {iopath_Amult26_Cmult42} {iopath_Amult26_Cmult43} {iopath_Amult26_Cmult44} {iopath_Amult26_Cmult45} {iopath_Amult26_Cmult46} {iopath_Amult26_Cmult47} {iopath_Amult26_Cmult48} {iopath_Amult26_Cmult49} {iopath_Amult26_Cmult50} {iopath_Amult26_Cmult51} {iopath_Amult26_Cmult52} {iopath_Amult26_Cmult53} {iopath_Amult26_Cmult54} {iopath_Amult26_Cmult55} {iopath_Amult26_Cmult56} {iopath_Amult26_Cmult57} {iopath_Amult26_Cmult58} {iopath_Amult26_Cmult59} {iopath_Amult26_Cmult60} {iopath_Amult26_Cmult61} {iopath_Amult26_Cmult62} {iopath_Amult26_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult27_Cmult27} {iopath_Amult27_Cmult28} {iopath_Amult27_Cmult29} {iopath_Amult27_Cmult30} {iopath_Amult27_Cmult31} {iopath_Amult27_Cmult32} {iopath_Amult27_Cmult33} {iopath_Amult27_Cmult34} {iopath_Amult27_Cmult35} {iopath_Amult27_Cmult36} {iopath_Amult27_Cmult37} {iopath_Amult27_Cmult38} {iopath_Amult27_Cmult39} {iopath_Amult27_Cmult40} {iopath_Amult27_Cmult41} {iopath_Amult27_Cmult42} {iopath_Amult27_Cmult43} {iopath_Amult27_Cmult44} {iopath_Amult27_Cmult45} {iopath_Amult27_Cmult46} {iopath_Amult27_Cmult47} {iopath_Amult27_Cmult48} {iopath_Amult27_Cmult49} {iopath_Amult27_Cmult50} {iopath_Amult27_Cmult51} {iopath_Amult27_Cmult52} {iopath_Amult27_Cmult53} {iopath_Amult27_Cmult54} {iopath_Amult27_Cmult55} {iopath_Amult27_Cmult56} {iopath_Amult27_Cmult57} {iopath_Amult27_Cmult58} {iopath_Amult27_Cmult59} {iopath_Amult27_Cmult60} {iopath_Amult27_Cmult61} {iopath_Amult27_Cmult62} {iopath_Amult27_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult28_Cmult28} {iopath_Amult28_Cmult29} {iopath_Amult28_Cmult30} {iopath_Amult28_Cmult31} {iopath_Amult28_Cmult32} {iopath_Amult28_Cmult33} {iopath_Amult28_Cmult34} {iopath_Amult28_Cmult35} {iopath_Amult28_Cmult36} {iopath_Amult28_Cmult37} {iopath_Amult28_Cmult38} {iopath_Amult28_Cmult39} {iopath_Amult28_Cmult40} {iopath_Amult28_Cmult41} {iopath_Amult28_Cmult42} {iopath_Amult28_Cmult43} {iopath_Amult28_Cmult44} {iopath_Amult28_Cmult45} {iopath_Amult28_Cmult46} {iopath_Amult28_Cmult47} {iopath_Amult28_Cmult48} {iopath_Amult28_Cmult49} {iopath_Amult28_Cmult50} {iopath_Amult28_Cmult51} {iopath_Amult28_Cmult52} {iopath_Amult28_Cmult53} {iopath_Amult28_Cmult54} {iopath_Amult28_Cmult55} {iopath_Amult28_Cmult56} {iopath_Amult28_Cmult57} {iopath_Amult28_Cmult58} {iopath_Amult28_Cmult59} {iopath_Amult28_Cmult60} {iopath_Amult28_Cmult61} {iopath_Amult28_Cmult62} {iopath_Amult28_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult29_Cmult29} {iopath_Amult29_Cmult30} {iopath_Amult29_Cmult31} {iopath_Amult29_Cmult32} {iopath_Amult29_Cmult33} {iopath_Amult29_Cmult34} {iopath_Amult29_Cmult35} {iopath_Amult29_Cmult36} {iopath_Amult29_Cmult37} {iopath_Amult29_Cmult38} {iopath_Amult29_Cmult39} {iopath_Amult29_Cmult40} {iopath_Amult29_Cmult41} {iopath_Amult29_Cmult42} {iopath_Amult29_Cmult43} {iopath_Amult29_Cmult44} {iopath_Amult29_Cmult45} {iopath_Amult29_Cmult46} {iopath_Amult29_Cmult47} {iopath_Amult29_Cmult48} {iopath_Amult29_Cmult49} {iopath_Amult29_Cmult50} {iopath_Amult29_Cmult51} {iopath_Amult29_Cmult52} {iopath_Amult29_Cmult53} {iopath_Amult29_Cmult54} {iopath_Amult29_Cmult55} {iopath_Amult29_Cmult56} {iopath_Amult29_Cmult57} {iopath_Amult29_Cmult58} {iopath_Amult29_Cmult59} {iopath_Amult29_Cmult60} {iopath_Amult29_Cmult61} {iopath_Amult29_Cmult62} {iopath_Amult29_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult30_Cmult30} {iopath_Amult30_Cmult31} {iopath_Amult30_Cmult32} {iopath_Amult30_Cmult33} {iopath_Amult30_Cmult34} {iopath_Amult30_Cmult35} {iopath_Amult30_Cmult36} {iopath_Amult30_Cmult37} {iopath_Amult30_Cmult38} {iopath_Amult30_Cmult39} {iopath_Amult30_Cmult40} {iopath_Amult30_Cmult41} {iopath_Amult30_Cmult42} {iopath_Amult30_Cmult43} {iopath_Amult30_Cmult44} {iopath_Amult30_Cmult45} {iopath_Amult30_Cmult46} {iopath_Amult30_Cmult47} {iopath_Amult30_Cmult48} {iopath_Amult30_Cmult49} {iopath_Amult30_Cmult50} {iopath_Amult30_Cmult51} {iopath_Amult30_Cmult52} {iopath_Amult30_Cmult53} {iopath_Amult30_Cmult54} {iopath_Amult30_Cmult55} {iopath_Amult30_Cmult56} {iopath_Amult30_Cmult57} {iopath_Amult30_Cmult58} {iopath_Amult30_Cmult59} {iopath_Amult30_Cmult60} {iopath_Amult30_Cmult61} {iopath_Amult30_Cmult62} {iopath_Amult30_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult31_Cmult31} {iopath_Amult31_Cmult32} {iopath_Amult31_Cmult33} {iopath_Amult31_Cmult34} {iopath_Amult31_Cmult35} {iopath_Amult31_Cmult36} {iopath_Amult31_Cmult37} {iopath_Amult31_Cmult38} {iopath_Amult31_Cmult39} {iopath_Amult31_Cmult40} {iopath_Amult31_Cmult41} {iopath_Amult31_Cmult42} {iopath_Amult31_Cmult43} {iopath_Amult31_Cmult44} {iopath_Amult31_Cmult45} {iopath_Amult31_Cmult46} {iopath_Amult31_Cmult47} {iopath_Amult31_Cmult48} {iopath_Amult31_Cmult49} {iopath_Amult31_Cmult50} {iopath_Amult31_Cmult51} {iopath_Amult31_Cmult52} {iopath_Amult31_Cmult53} {iopath_Amult31_Cmult54} {iopath_Amult31_Cmult55} {iopath_Amult31_Cmult56} {iopath_Amult31_Cmult57} {iopath_Amult31_Cmult58} {iopath_Amult31_Cmult59} {iopath_Amult31_Cmult60} {iopath_Amult31_Cmult61} {iopath_Amult31_Cmult62} {iopath_Amult31_Cmult63} "*)
	(* DELAY_MATRIX_Bmult="{iopath_Amult0_Cmult0} {iopath_Amult0_Cmult1} {iopath_Amult0_Cmult2} {iopath_Amult0_Cmult3} {iopath_Amult0_Cmult4} {iopath_Amult0_Cmult5} {iopath_Amult0_Cmult6} {iopath_Amult0_Cmult7} {iopath_Amult0_Cmult8} {iopath_Amult0_Cmult9} {iopath_Amult0_Cmult10} {iopath_Amult0_Cmult11} {iopath_Amult0_Cmult12} {iopath_Amult0_Cmult13} {iopath_Amult0_Cmult14} {iopath_Amult0_Cmult15} {iopath_Amult0_Cmult16} {iopath_Amult0_Cmult17} {iopath_Amult0_Cmult18} {iopath_Amult0_Cmult19} {iopath_Amult0_Cmult20} {iopath_Amult0_Cmult21} {iopath_Amult0_Cmult22} {iopath_Amult0_Cmult23} {iopath_Amult0_Cmult24} {iopath_Amult0_Cmult25} {iopath_Amult0_Cmult26} {iopath_Amult0_Cmult27} {iopath_Amult0_Cmult28} {iopath_Amult0_Cmult29} {iopath_Amult0_Cmult30} {iopath_Amult0_Cmult31} {iopath_Amult0_Cmult32} {iopath_Amult0_Cmult33} {iopath_Amult0_Cmult34} {iopath_Amult0_Cmult35} {iopath_Amult0_Cmult36} {iopath_Amult0_Cmult37} {iopath_Amult0_Cmult38} {iopath_Amult0_Cmult39} {iopath_Amult0_Cmult40} {iopath_Amult0_Cmult41} {iopath_Amult0_Cmult42} {iopath_Amult0_Cmult43} {iopath_Amult0_Cmult44} {iopath_Amult0_Cmult45} {iopath_Amult0_Cmult46} {iopath_Amult0_Cmult47} {iopath_Amult0_Cmult48} {iopath_Amult0_Cmult49} {iopath_Amult0_Cmult50} {iopath_Amult0_Cmult51} {iopath_Amult0_Cmult52} {iopath_Amult0_Cmult53} {iopath_Amult0_Cmult54} {iopath_Amult0_Cmult55} {iopath_Amult0_Cmult56} {iopath_Amult0_Cmult57} {iopath_Amult0_Cmult58} {iopath_Amult0_Cmult59} {iopath_Amult0_Cmult60} {iopath_Amult0_Cmult61} {iopath_Amult0_Cmult62} {iopath_Amult0_Cmult63} 0 {iopath_Amult1_Cmult1} {iopath_Amult1_Cmult2} {iopath_Amult1_Cmult3} {iopath_Amult1_Cmult4} {iopath_Amult1_Cmult5} {iopath_Amult1_Cmult6} {iopath_Amult1_Cmult7} {iopath_Amult1_Cmult8} {iopath_Amult1_Cmult9} {iopath_Amult1_Cmult10} {iopath_Amult1_Cmult11} {iopath_Amult1_Cmult12} {iopath_Amult1_Cmult13} {iopath_Amult1_Cmult14} {iopath_Amult1_Cmult15} {iopath_Amult1_Cmult16} {iopath_Amult1_Cmult17} {iopath_Amult1_Cmult18} {iopath_Amult1_Cmult19} {iopath_Amult1_Cmult20} {iopath_Amult1_Cmult21} {iopath_Amult1_Cmult22} {iopath_Amult1_Cmult23} {iopath_Amult1_Cmult24} {iopath_Amult1_Cmult25} {iopath_Amult1_Cmult26} {iopath_Amult1_Cmult27} {iopath_Amult1_Cmult28} {iopath_Amult1_Cmult29} {iopath_Amult1_Cmult30} {iopath_Amult1_Cmult31} {iopath_Amult1_Cmult32} {iopath_Amult1_Cmult33} {iopath_Amult1_Cmult34} {iopath_Amult1_Cmult35} {iopath_Amult1_Cmult36} {iopath_Amult1_Cmult37} {iopath_Amult1_Cmult38} {iopath_Amult1_Cmult39} {iopath_Amult1_Cmult40} {iopath_Amult1_Cmult41} {iopath_Amult1_Cmult42} {iopath_Amult1_Cmult43} {iopath_Amult1_Cmult44} {iopath_Amult1_Cmult45} {iopath_Amult1_Cmult46} {iopath_Amult1_Cmult47} {iopath_Amult1_Cmult48} {iopath_Amult1_Cmult49} {iopath_Amult1_Cmult50} {iopath_Amult1_Cmult51} {iopath_Amult1_Cmult52} {iopath_Amult1_Cmult53} {iopath_Amult1_Cmult54} {iopath_Amult1_Cmult55} {iopath_Amult1_Cmult56} {iopath_Amult1_Cmult57} {iopath_Amult1_Cmult58} {iopath_Amult1_Cmult59} {iopath_Amult1_Cmult60} {iopath_Amult1_Cmult61} {iopath_Amult1_Cmult62} {iopath_Amult1_Cmult63} 0 0 {iopath_Amult2_Cmult2} {iopath_Amult2_Cmult3} {iopath_Amult2_Cmult4} {iopath_Amult2_Cmult5} {iopath_Amult2_Cmult6} {iopath_Amult2_Cmult7} {iopath_Amult2_Cmult8} {iopath_Amult2_Cmult9} {iopath_Amult2_Cmult10} {iopath_Amult2_Cmult11} {iopath_Amult2_Cmult12} {iopath_Amult2_Cmult13} {iopath_Amult2_Cmult14} {iopath_Amult2_Cmult15} {iopath_Amult2_Cmult16} {iopath_Amult2_Cmult17} {iopath_Amult2_Cmult18} {iopath_Amult2_Cmult19} {iopath_Amult2_Cmult20} {iopath_Amult2_Cmult21} {iopath_Amult2_Cmult22} {iopath_Amult2_Cmult23} {iopath_Amult2_Cmult24} {iopath_Amult2_Cmult25} {iopath_Amult2_Cmult26} {iopath_Amult2_Cmult27} {iopath_Amult2_Cmult28} {iopath_Amult2_Cmult29} {iopath_Amult2_Cmult30} {iopath_Amult2_Cmult31} {iopath_Amult2_Cmult32} {iopath_Amult2_Cmult33} {iopath_Amult2_Cmult34} {iopath_Amult2_Cmult35} {iopath_Amult2_Cmult36} {iopath_Amult2_Cmult37} {iopath_Amult2_Cmult38} {iopath_Amult2_Cmult39} {iopath_Amult2_Cmult40} {iopath_Amult2_Cmult41} {iopath_Amult2_Cmult42} {iopath_Amult2_Cmult43} {iopath_Amult2_Cmult44} {iopath_Amult2_Cmult45} {iopath_Amult2_Cmult46} {iopath_Amult2_Cmult47} {iopath_Amult2_Cmult48} {iopath_Amult2_Cmult49} {iopath_Amult2_Cmult50} {iopath_Amult2_Cmult51} {iopath_Amult2_Cmult52} {iopath_Amult2_Cmult53} {iopath_Amult2_Cmult54} {iopath_Amult2_Cmult55} {iopath_Amult2_Cmult56} {iopath_Amult2_Cmult57} {iopath_Amult2_Cmult58} {iopath_Amult2_Cmult59} {iopath_Amult2_Cmult60} {iopath_Amult2_Cmult61} {iopath_Amult2_Cmult62} {iopath_Amult2_Cmult63} 0 0 0 {iopath_Amult3_Cmult3} {iopath_Amult3_Cmult4} {iopath_Amult3_Cmult5} {iopath_Amult3_Cmult6} {iopath_Amult3_Cmult7} {iopath_Amult3_Cmult8} {iopath_Amult3_Cmult9} {iopath_Amult3_Cmult10} {iopath_Amult3_Cmult11} {iopath_Amult3_Cmult12} {iopath_Amult3_Cmult13} {iopath_Amult3_Cmult14} {iopath_Amult3_Cmult15} {iopath_Amult3_Cmult16} {iopath_Amult3_Cmult17} {iopath_Amult3_Cmult18} {iopath_Amult3_Cmult19} {iopath_Amult3_Cmult20} {iopath_Amult3_Cmult21} {iopath_Amult3_Cmult22} {iopath_Amult3_Cmult23} {iopath_Amult3_Cmult24} {iopath_Amult3_Cmult25} {iopath_Amult3_Cmult26} {iopath_Amult3_Cmult27} {iopath_Amult3_Cmult28} {iopath_Amult3_Cmult29} {iopath_Amult3_Cmult30} {iopath_Amult3_Cmult31} {iopath_Amult3_Cmult32} {iopath_Amult3_Cmult33} {iopath_Amult3_Cmult34} {iopath_Amult3_Cmult35} {iopath_Amult3_Cmult36} {iopath_Amult3_Cmult37} {iopath_Amult3_Cmult38} {iopath_Amult3_Cmult39} {iopath_Amult3_Cmult40} {iopath_Amult3_Cmult41} {iopath_Amult3_Cmult42} {iopath_Amult3_Cmult43} {iopath_Amult3_Cmult44} {iopath_Amult3_Cmult45} {iopath_Amult3_Cmult46} {iopath_Amult3_Cmult47} {iopath_Amult3_Cmult48} {iopath_Amult3_Cmult49} {iopath_Amult3_Cmult50} {iopath_Amult3_Cmult51} {iopath_Amult3_Cmult52} {iopath_Amult3_Cmult53} {iopath_Amult3_Cmult54} {iopath_Amult3_Cmult55} {iopath_Amult3_Cmult56} {iopath_Amult3_Cmult57} {iopath_Amult3_Cmult58} {iopath_Amult3_Cmult59} {iopath_Amult3_Cmult60} {iopath_Amult3_Cmult61} {iopath_Amult3_Cmult62} {iopath_Amult3_Cmult63} 0 0 0 0 {iopath_Amult4_Cmult4} {iopath_Amult4_Cmult5} {iopath_Amult4_Cmult6} {iopath_Amult4_Cmult7} {iopath_Amult4_Cmult8} {iopath_Amult4_Cmult9} {iopath_Amult4_Cmult10} {iopath_Amult4_Cmult11} {iopath_Amult4_Cmult12} {iopath_Amult4_Cmult13} {iopath_Amult4_Cmult14} {iopath_Amult4_Cmult15} {iopath_Amult4_Cmult16} {iopath_Amult4_Cmult17} {iopath_Amult4_Cmult18} {iopath_Amult4_Cmult19} {iopath_Amult4_Cmult20} {iopath_Amult4_Cmult21} {iopath_Amult4_Cmult22} {iopath_Amult4_Cmult23} {iopath_Amult4_Cmult24} {iopath_Amult4_Cmult25} {iopath_Amult4_Cmult26} {iopath_Amult4_Cmult27} {iopath_Amult4_Cmult28} {iopath_Amult4_Cmult29} {iopath_Amult4_Cmult30} {iopath_Amult4_Cmult31} {iopath_Amult4_Cmult32} {iopath_Amult4_Cmult33} {iopath_Amult4_Cmult34} {iopath_Amult4_Cmult35} {iopath_Amult4_Cmult36} {iopath_Amult4_Cmult37} {iopath_Amult4_Cmult38} {iopath_Amult4_Cmult39} {iopath_Amult4_Cmult40} {iopath_Amult4_Cmult41} {iopath_Amult4_Cmult42} {iopath_Amult4_Cmult43} {iopath_Amult4_Cmult44} {iopath_Amult4_Cmult45} {iopath_Amult4_Cmult46} {iopath_Amult4_Cmult47} {iopath_Amult4_Cmult48} {iopath_Amult4_Cmult49} {iopath_Amult4_Cmult50} {iopath_Amult4_Cmult51} {iopath_Amult4_Cmult52} {iopath_Amult4_Cmult53} {iopath_Amult4_Cmult54} {iopath_Amult4_Cmult55} {iopath_Amult4_Cmult56} {iopath_Amult4_Cmult57} {iopath_Amult4_Cmult58} {iopath_Amult4_Cmult59} {iopath_Amult4_Cmult60} {iopath_Amult4_Cmult61} {iopath_Amult4_Cmult62} {iopath_Amult4_Cmult63} 0 0 0 0 0 {iopath_Amult5_Cmult5} {iopath_Amult5_Cmult6} {iopath_Amult5_Cmult7} {iopath_Amult5_Cmult8} {iopath_Amult5_Cmult9} {iopath_Amult5_Cmult10} {iopath_Amult5_Cmult11} {iopath_Amult5_Cmult12} {iopath_Amult5_Cmult13} {iopath_Amult5_Cmult14} {iopath_Amult5_Cmult15} {iopath_Amult5_Cmult16} {iopath_Amult5_Cmult17} {iopath_Amult5_Cmult18} {iopath_Amult5_Cmult19} {iopath_Amult5_Cmult20} {iopath_Amult5_Cmult21} {iopath_Amult5_Cmult22} {iopath_Amult5_Cmult23} {iopath_Amult5_Cmult24} {iopath_Amult5_Cmult25} {iopath_Amult5_Cmult26} {iopath_Amult5_Cmult27} {iopath_Amult5_Cmult28} {iopath_Amult5_Cmult29} {iopath_Amult5_Cmult30} {iopath_Amult5_Cmult31} {iopath_Amult5_Cmult32} {iopath_Amult5_Cmult33} {iopath_Amult5_Cmult34} {iopath_Amult5_Cmult35} {iopath_Amult5_Cmult36} {iopath_Amult5_Cmult37} {iopath_Amult5_Cmult38} {iopath_Amult5_Cmult39} {iopath_Amult5_Cmult40} {iopath_Amult5_Cmult41} {iopath_Amult5_Cmult42} {iopath_Amult5_Cmult43} {iopath_Amult5_Cmult44} {iopath_Amult5_Cmult45} {iopath_Amult5_Cmult46} {iopath_Amult5_Cmult47} {iopath_Amult5_Cmult48} {iopath_Amult5_Cmult49} {iopath_Amult5_Cmult50} {iopath_Amult5_Cmult51} {iopath_Amult5_Cmult52} {iopath_Amult5_Cmult53} {iopath_Amult5_Cmult54} {iopath_Amult5_Cmult55} {iopath_Amult5_Cmult56} {iopath_Amult5_Cmult57} {iopath_Amult5_Cmult58} {iopath_Amult5_Cmult59} {iopath_Amult5_Cmult60} {iopath_Amult5_Cmult61} {iopath_Amult5_Cmult62} {iopath_Amult5_Cmult63} 0 0 0 0 0 0 {iopath_Amult6_Cmult6} {iopath_Amult6_Cmult7} {iopath_Amult6_Cmult8} {iopath_Amult6_Cmult9} {iopath_Amult6_Cmult10} {iopath_Amult6_Cmult11} {iopath_Amult6_Cmult12} {iopath_Amult6_Cmult13} {iopath_Amult6_Cmult14} {iopath_Amult6_Cmult15} {iopath_Amult6_Cmult16} {iopath_Amult6_Cmult17} {iopath_Amult6_Cmult18} {iopath_Amult6_Cmult19} {iopath_Amult6_Cmult20} {iopath_Amult6_Cmult21} {iopath_Amult6_Cmult22} {iopath_Amult6_Cmult23} {iopath_Amult6_Cmult24} {iopath_Amult6_Cmult25} {iopath_Amult6_Cmult26} {iopath_Amult6_Cmult27} {iopath_Amult6_Cmult28} {iopath_Amult6_Cmult29} {iopath_Amult6_Cmult30} {iopath_Amult6_Cmult31} {iopath_Amult6_Cmult32} {iopath_Amult6_Cmult33} {iopath_Amult6_Cmult34} {iopath_Amult6_Cmult35} {iopath_Amult6_Cmult36} {iopath_Amult6_Cmult37} {iopath_Amult6_Cmult38} {iopath_Amult6_Cmult39} {iopath_Amult6_Cmult40} {iopath_Amult6_Cmult41} {iopath_Amult6_Cmult42} {iopath_Amult6_Cmult43} {iopath_Amult6_Cmult44} {iopath_Amult6_Cmult45} {iopath_Amult6_Cmult46} {iopath_Amult6_Cmult47} {iopath_Amult6_Cmult48} {iopath_Amult6_Cmult49} {iopath_Amult6_Cmult50} {iopath_Amult6_Cmult51} {iopath_Amult6_Cmult52} {iopath_Amult6_Cmult53} {iopath_Amult6_Cmult54} {iopath_Amult6_Cmult55} {iopath_Amult6_Cmult56} {iopath_Amult6_Cmult57} {iopath_Amult6_Cmult58} {iopath_Amult6_Cmult59} {iopath_Amult6_Cmult60} {iopath_Amult6_Cmult61} {iopath_Amult6_Cmult62} {iopath_Amult6_Cmult63} 0 0 0 0 0 0 0 {iopath_Amult7_Cmult7} {iopath_Amult7_Cmult8} {iopath_Amult7_Cmult9} {iopath_Amult7_Cmult10} {iopath_Amult7_Cmult11} {iopath_Amult7_Cmult12} {iopath_Amult7_Cmult13} {iopath_Amult7_Cmult14} {iopath_Amult7_Cmult15} {iopath_Amult7_Cmult16} {iopath_Amult7_Cmult17} {iopath_Amult7_Cmult18} {iopath_Amult7_Cmult19} {iopath_Amult7_Cmult20} {iopath_Amult7_Cmult21} {iopath_Amult7_Cmult22} {iopath_Amult7_Cmult23} {iopath_Amult7_Cmult24} {iopath_Amult7_Cmult25} {iopath_Amult7_Cmult26} {iopath_Amult7_Cmult27} {iopath_Amult7_Cmult28} {iopath_Amult7_Cmult29} {iopath_Amult7_Cmult30} {iopath_Amult7_Cmult31} {iopath_Amult7_Cmult32} {iopath_Amult7_Cmult33} {iopath_Amult7_Cmult34} {iopath_Amult7_Cmult35} {iopath_Amult7_Cmult36} {iopath_Amult7_Cmult37} {iopath_Amult7_Cmult38} {iopath_Amult7_Cmult39} {iopath_Amult7_Cmult40} {iopath_Amult7_Cmult41} {iopath_Amult7_Cmult42} {iopath_Amult7_Cmult43} {iopath_Amult7_Cmult44} {iopath_Amult7_Cmult45} {iopath_Amult7_Cmult46} {iopath_Amult7_Cmult47} {iopath_Amult7_Cmult48} {iopath_Amult7_Cmult49} {iopath_Amult7_Cmult50} {iopath_Amult7_Cmult51} {iopath_Amult7_Cmult52} {iopath_Amult7_Cmult53} {iopath_Amult7_Cmult54} {iopath_Amult7_Cmult55} {iopath_Amult7_Cmult56} {iopath_Amult7_Cmult57} {iopath_Amult7_Cmult58} {iopath_Amult7_Cmult59} {iopath_Amult7_Cmult60} {iopath_Amult7_Cmult61} {iopath_Amult7_Cmult62} {iopath_Amult7_Cmult63} 0 0 0 0 0 0 0 0 {iopath_Amult8_Cmult8} {iopath_Amult8_Cmult9} {iopath_Amult8_Cmult10} {iopath_Amult8_Cmult11} {iopath_Amult8_Cmult12} {iopath_Amult8_Cmult13} {iopath_Amult8_Cmult14} {iopath_Amult8_Cmult15} {iopath_Amult8_Cmult16} {iopath_Amult8_Cmult17} {iopath_Amult8_Cmult18} {iopath_Amult8_Cmult19} {iopath_Amult8_Cmult20} {iopath_Amult8_Cmult21} {iopath_Amult8_Cmult22} {iopath_Amult8_Cmult23} {iopath_Amult8_Cmult24} {iopath_Amult8_Cmult25} {iopath_Amult8_Cmult26} {iopath_Amult8_Cmult27} {iopath_Amult8_Cmult28} {iopath_Amult8_Cmult29} {iopath_Amult8_Cmult30} {iopath_Amult8_Cmult31} {iopath_Amult8_Cmult32} {iopath_Amult8_Cmult33} {iopath_Amult8_Cmult34} {iopath_Amult8_Cmult35} {iopath_Amult8_Cmult36} {iopath_Amult8_Cmult37} {iopath_Amult8_Cmult38} {iopath_Amult8_Cmult39} {iopath_Amult8_Cmult40} {iopath_Amult8_Cmult41} {iopath_Amult8_Cmult42} {iopath_Amult8_Cmult43} {iopath_Amult8_Cmult44} {iopath_Amult8_Cmult45} {iopath_Amult8_Cmult46} {iopath_Amult8_Cmult47} {iopath_Amult8_Cmult48} {iopath_Amult8_Cmult49} {iopath_Amult8_Cmult50} {iopath_Amult8_Cmult51} {iopath_Amult8_Cmult52} {iopath_Amult8_Cmult53} {iopath_Amult8_Cmult54} {iopath_Amult8_Cmult55} {iopath_Amult8_Cmult56} {iopath_Amult8_Cmult57} {iopath_Amult8_Cmult58} {iopath_Amult8_Cmult59} {iopath_Amult8_Cmult60} {iopath_Amult8_Cmult61} {iopath_Amult8_Cmult62} {iopath_Amult8_Cmult63} 0 0 0 0 0 0 0 0 0 {iopath_Amult9_Cmult9} {iopath_Amult9_Cmult10} {iopath_Amult9_Cmult11} {iopath_Amult9_Cmult12} {iopath_Amult9_Cmult13} {iopath_Amult9_Cmult14} {iopath_Amult9_Cmult15} {iopath_Amult9_Cmult16} {iopath_Amult9_Cmult17} {iopath_Amult9_Cmult18} {iopath_Amult9_Cmult19} {iopath_Amult9_Cmult20} {iopath_Amult9_Cmult21} {iopath_Amult9_Cmult22} {iopath_Amult9_Cmult23} {iopath_Amult9_Cmult24} {iopath_Amult9_Cmult25} {iopath_Amult9_Cmult26} {iopath_Amult9_Cmult27} {iopath_Amult9_Cmult28} {iopath_Amult9_Cmult29} {iopath_Amult9_Cmult30} {iopath_Amult9_Cmult31} {iopath_Amult9_Cmult32} {iopath_Amult9_Cmult33} {iopath_Amult9_Cmult34} {iopath_Amult9_Cmult35} {iopath_Amult9_Cmult36} {iopath_Amult9_Cmult37} {iopath_Amult9_Cmult38} {iopath_Amult9_Cmult39} {iopath_Amult9_Cmult40} {iopath_Amult9_Cmult41} {iopath_Amult9_Cmult42} {iopath_Amult9_Cmult43} {iopath_Amult9_Cmult44} {iopath_Amult9_Cmult45} {iopath_Amult9_Cmult46} {iopath_Amult9_Cmult47} {iopath_Amult9_Cmult48} {iopath_Amult9_Cmult49} {iopath_Amult9_Cmult50} {iopath_Amult9_Cmult51} {iopath_Amult9_Cmult52} {iopath_Amult9_Cmult53} {iopath_Amult9_Cmult54} {iopath_Amult9_Cmult55} {iopath_Amult9_Cmult56} {iopath_Amult9_Cmult57} {iopath_Amult9_Cmult58} {iopath_Amult9_Cmult59} {iopath_Amult9_Cmult60} {iopath_Amult9_Cmult61} {iopath_Amult9_Cmult62} {iopath_Amult9_Cmult63} 0 0 0 0 0 0 0 0 0 0 {iopath_Amult10_Cmult10} {iopath_Amult10_Cmult11} {iopath_Amult10_Cmult12} {iopath_Amult10_Cmult13} {iopath_Amult10_Cmult14} {iopath_Amult10_Cmult15} {iopath_Amult10_Cmult16} {iopath_Amult10_Cmult17} {iopath_Amult10_Cmult18} {iopath_Amult10_Cmult19} {iopath_Amult10_Cmult20} {iopath_Amult10_Cmult21} {iopath_Amult10_Cmult22} {iopath_Amult10_Cmult23} {iopath_Amult10_Cmult24} {iopath_Amult10_Cmult25} {iopath_Amult10_Cmult26} {iopath_Amult10_Cmult27} {iopath_Amult10_Cmult28} {iopath_Amult10_Cmult29} {iopath_Amult10_Cmult30} {iopath_Amult10_Cmult31} {iopath_Amult10_Cmult32} {iopath_Amult10_Cmult33} {iopath_Amult10_Cmult34} {iopath_Amult10_Cmult35} {iopath_Amult10_Cmult36} {iopath_Amult10_Cmult37} {iopath_Amult10_Cmult38} {iopath_Amult10_Cmult39} {iopath_Amult10_Cmult40} {iopath_Amult10_Cmult41} {iopath_Amult10_Cmult42} {iopath_Amult10_Cmult43} {iopath_Amult10_Cmult44} {iopath_Amult10_Cmult45} {iopath_Amult10_Cmult46} {iopath_Amult10_Cmult47} {iopath_Amult10_Cmult48} {iopath_Amult10_Cmult49} {iopath_Amult10_Cmult50} {iopath_Amult10_Cmult51} {iopath_Amult10_Cmult52} {iopath_Amult10_Cmult53} {iopath_Amult10_Cmult54} {iopath_Amult10_Cmult55} {iopath_Amult10_Cmult56} {iopath_Amult10_Cmult57} {iopath_Amult10_Cmult58} {iopath_Amult10_Cmult59} {iopath_Amult10_Cmult60} {iopath_Amult10_Cmult61} {iopath_Amult10_Cmult62} {iopath_Amult10_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult11_Cmult11} {iopath_Amult11_Cmult12} {iopath_Amult11_Cmult13} {iopath_Amult11_Cmult14} {iopath_Amult11_Cmult15} {iopath_Amult11_Cmult16} {iopath_Amult11_Cmult17} {iopath_Amult11_Cmult18} {iopath_Amult11_Cmult19} {iopath_Amult11_Cmult20} {iopath_Amult11_Cmult21} {iopath_Amult11_Cmult22} {iopath_Amult11_Cmult23} {iopath_Amult11_Cmult24} {iopath_Amult11_Cmult25} {iopath_Amult11_Cmult26} {iopath_Amult11_Cmult27} {iopath_Amult11_Cmult28} {iopath_Amult11_Cmult29} {iopath_Amult11_Cmult30} {iopath_Amult11_Cmult31} {iopath_Amult11_Cmult32} {iopath_Amult11_Cmult33} {iopath_Amult11_Cmult34} {iopath_Amult11_Cmult35} {iopath_Amult11_Cmult36} {iopath_Amult11_Cmult37} {iopath_Amult11_Cmult38} {iopath_Amult11_Cmult39} {iopath_Amult11_Cmult40} {iopath_Amult11_Cmult41} {iopath_Amult11_Cmult42} {iopath_Amult11_Cmult43} {iopath_Amult11_Cmult44} {iopath_Amult11_Cmult45} {iopath_Amult11_Cmult46} {iopath_Amult11_Cmult47} {iopath_Amult11_Cmult48} {iopath_Amult11_Cmult49} {iopath_Amult11_Cmult50} {iopath_Amult11_Cmult51} {iopath_Amult11_Cmult52} {iopath_Amult11_Cmult53} {iopath_Amult11_Cmult54} {iopath_Amult11_Cmult55} {iopath_Amult11_Cmult56} {iopath_Amult11_Cmult57} {iopath_Amult11_Cmult58} {iopath_Amult11_Cmult59} {iopath_Amult11_Cmult60} {iopath_Amult11_Cmult61} {iopath_Amult11_Cmult62} {iopath_Amult11_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult12_Cmult12} {iopath_Amult12_Cmult13} {iopath_Amult12_Cmult14} {iopath_Amult12_Cmult15} {iopath_Amult12_Cmult16} {iopath_Amult12_Cmult17} {iopath_Amult12_Cmult18} {iopath_Amult12_Cmult19} {iopath_Amult12_Cmult20} {iopath_Amult12_Cmult21} {iopath_Amult12_Cmult22} {iopath_Amult12_Cmult23} {iopath_Amult12_Cmult24} {iopath_Amult12_Cmult25} {iopath_Amult12_Cmult26} {iopath_Amult12_Cmult27} {iopath_Amult12_Cmult28} {iopath_Amult12_Cmult29} {iopath_Amult12_Cmult30} {iopath_Amult12_Cmult31} {iopath_Amult12_Cmult32} {iopath_Amult12_Cmult33} {iopath_Amult12_Cmult34} {iopath_Amult12_Cmult35} {iopath_Amult12_Cmult36} {iopath_Amult12_Cmult37} {iopath_Amult12_Cmult38} {iopath_Amult12_Cmult39} {iopath_Amult12_Cmult40} {iopath_Amult12_Cmult41} {iopath_Amult12_Cmult42} {iopath_Amult12_Cmult43} {iopath_Amult12_Cmult44} {iopath_Amult12_Cmult45} {iopath_Amult12_Cmult46} {iopath_Amult12_Cmult47} {iopath_Amult12_Cmult48} {iopath_Amult12_Cmult49} {iopath_Amult12_Cmult50} {iopath_Amult12_Cmult51} {iopath_Amult12_Cmult52} {iopath_Amult12_Cmult53} {iopath_Amult12_Cmult54} {iopath_Amult12_Cmult55} {iopath_Amult12_Cmult56} {iopath_Amult12_Cmult57} {iopath_Amult12_Cmult58} {iopath_Amult12_Cmult59} {iopath_Amult12_Cmult60} {iopath_Amult12_Cmult61} {iopath_Amult12_Cmult62} {iopath_Amult12_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult13_Cmult13} {iopath_Amult13_Cmult14} {iopath_Amult13_Cmult15} {iopath_Amult13_Cmult16} {iopath_Amult13_Cmult17} {iopath_Amult13_Cmult18} {iopath_Amult13_Cmult19} {iopath_Amult13_Cmult20} {iopath_Amult13_Cmult21} {iopath_Amult13_Cmult22} {iopath_Amult13_Cmult23} {iopath_Amult13_Cmult24} {iopath_Amult13_Cmult25} {iopath_Amult13_Cmult26} {iopath_Amult13_Cmult27} {iopath_Amult13_Cmult28} {iopath_Amult13_Cmult29} {iopath_Amult13_Cmult30} {iopath_Amult13_Cmult31} {iopath_Amult13_Cmult32} {iopath_Amult13_Cmult33} {iopath_Amult13_Cmult34} {iopath_Amult13_Cmult35} {iopath_Amult13_Cmult36} {iopath_Amult13_Cmult37} {iopath_Amult13_Cmult38} {iopath_Amult13_Cmult39} {iopath_Amult13_Cmult40} {iopath_Amult13_Cmult41} {iopath_Amult13_Cmult42} {iopath_Amult13_Cmult43} {iopath_Amult13_Cmult44} {iopath_Amult13_Cmult45} {iopath_Amult13_Cmult46} {iopath_Amult13_Cmult47} {iopath_Amult13_Cmult48} {iopath_Amult13_Cmult49} {iopath_Amult13_Cmult50} {iopath_Amult13_Cmult51} {iopath_Amult13_Cmult52} {iopath_Amult13_Cmult53} {iopath_Amult13_Cmult54} {iopath_Amult13_Cmult55} {iopath_Amult13_Cmult56} {iopath_Amult13_Cmult57} {iopath_Amult13_Cmult58} {iopath_Amult13_Cmult59} {iopath_Amult13_Cmult60} {iopath_Amult13_Cmult61} {iopath_Amult13_Cmult62} {iopath_Amult13_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult14_Cmult14} {iopath_Amult14_Cmult15} {iopath_Amult14_Cmult16} {iopath_Amult14_Cmult17} {iopath_Amult14_Cmult18} {iopath_Amult14_Cmult19} {iopath_Amult14_Cmult20} {iopath_Amult14_Cmult21} {iopath_Amult14_Cmult22} {iopath_Amult14_Cmult23} {iopath_Amult14_Cmult24} {iopath_Amult14_Cmult25} {iopath_Amult14_Cmult26} {iopath_Amult14_Cmult27} {iopath_Amult14_Cmult28} {iopath_Amult14_Cmult29} {iopath_Amult14_Cmult30} {iopath_Amult14_Cmult31} {iopath_Amult14_Cmult32} {iopath_Amult14_Cmult33} {iopath_Amult14_Cmult34} {iopath_Amult14_Cmult35} {iopath_Amult14_Cmult36} {iopath_Amult14_Cmult37} {iopath_Amult14_Cmult38} {iopath_Amult14_Cmult39} {iopath_Amult14_Cmult40} {iopath_Amult14_Cmult41} {iopath_Amult14_Cmult42} {iopath_Amult14_Cmult43} {iopath_Amult14_Cmult44} {iopath_Amult14_Cmult45} {iopath_Amult14_Cmult46} {iopath_Amult14_Cmult47} {iopath_Amult14_Cmult48} {iopath_Amult14_Cmult49} {iopath_Amult14_Cmult50} {iopath_Amult14_Cmult51} {iopath_Amult14_Cmult52} {iopath_Amult14_Cmult53} {iopath_Amult14_Cmult54} {iopath_Amult14_Cmult55} {iopath_Amult14_Cmult56} {iopath_Amult14_Cmult57} {iopath_Amult14_Cmult58} {iopath_Amult14_Cmult59} {iopath_Amult14_Cmult60} {iopath_Amult14_Cmult61} {iopath_Amult14_Cmult62} {iopath_Amult14_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult15_Cmult15} {iopath_Amult15_Cmult16} {iopath_Amult15_Cmult17} {iopath_Amult15_Cmult18} {iopath_Amult15_Cmult19} {iopath_Amult15_Cmult20} {iopath_Amult15_Cmult21} {iopath_Amult15_Cmult22} {iopath_Amult15_Cmult23} {iopath_Amult15_Cmult24} {iopath_Amult15_Cmult25} {iopath_Amult15_Cmult26} {iopath_Amult15_Cmult27} {iopath_Amult15_Cmult28} {iopath_Amult15_Cmult29} {iopath_Amult15_Cmult30} {iopath_Amult15_Cmult31} {iopath_Amult15_Cmult32} {iopath_Amult15_Cmult33} {iopath_Amult15_Cmult34} {iopath_Amult15_Cmult35} {iopath_Amult15_Cmult36} {iopath_Amult15_Cmult37} {iopath_Amult15_Cmult38} {iopath_Amult15_Cmult39} {iopath_Amult15_Cmult40} {iopath_Amult15_Cmult41} {iopath_Amult15_Cmult42} {iopath_Amult15_Cmult43} {iopath_Amult15_Cmult44} {iopath_Amult15_Cmult45} {iopath_Amult15_Cmult46} {iopath_Amult15_Cmult47} {iopath_Amult15_Cmult48} {iopath_Amult15_Cmult49} {iopath_Amult15_Cmult50} {iopath_Amult15_Cmult51} {iopath_Amult15_Cmult52} {iopath_Amult15_Cmult53} {iopath_Amult15_Cmult54} {iopath_Amult15_Cmult55} {iopath_Amult15_Cmult56} {iopath_Amult15_Cmult57} {iopath_Amult15_Cmult58} {iopath_Amult15_Cmult59} {iopath_Amult15_Cmult60} {iopath_Amult15_Cmult61} {iopath_Amult15_Cmult62} {iopath_Amult15_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult16_Cmult16} {iopath_Amult16_Cmult17} {iopath_Amult16_Cmult18} {iopath_Amult16_Cmult19} {iopath_Amult16_Cmult20} {iopath_Amult16_Cmult21} {iopath_Amult16_Cmult22} {iopath_Amult16_Cmult23} {iopath_Amult16_Cmult24} {iopath_Amult16_Cmult25} {iopath_Amult16_Cmult26} {iopath_Amult16_Cmult27} {iopath_Amult16_Cmult28} {iopath_Amult16_Cmult29} {iopath_Amult16_Cmult30} {iopath_Amult16_Cmult31} {iopath_Amult16_Cmult32} {iopath_Amult16_Cmult33} {iopath_Amult16_Cmult34} {iopath_Amult16_Cmult35} {iopath_Amult16_Cmult36} {iopath_Amult16_Cmult37} {iopath_Amult16_Cmult38} {iopath_Amult16_Cmult39} {iopath_Amult16_Cmult40} {iopath_Amult16_Cmult41} {iopath_Amult16_Cmult42} {iopath_Amult16_Cmult43} {iopath_Amult16_Cmult44} {iopath_Amult16_Cmult45} {iopath_Amult16_Cmult46} {iopath_Amult16_Cmult47} {iopath_Amult16_Cmult48} {iopath_Amult16_Cmult49} {iopath_Amult16_Cmult50} {iopath_Amult16_Cmult51} {iopath_Amult16_Cmult52} {iopath_Amult16_Cmult53} {iopath_Amult16_Cmult54} {iopath_Amult16_Cmult55} {iopath_Amult16_Cmult56} {iopath_Amult16_Cmult57} {iopath_Amult16_Cmult58} {iopath_Amult16_Cmult59} {iopath_Amult16_Cmult60} {iopath_Amult16_Cmult61} {iopath_Amult16_Cmult62} {iopath_Amult16_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult17_Cmult17} {iopath_Amult17_Cmult18} {iopath_Amult17_Cmult19} {iopath_Amult17_Cmult20} {iopath_Amult17_Cmult21} {iopath_Amult17_Cmult22} {iopath_Amult17_Cmult23} {iopath_Amult17_Cmult24} {iopath_Amult17_Cmult25} {iopath_Amult17_Cmult26} {iopath_Amult17_Cmult27} {iopath_Amult17_Cmult28} {iopath_Amult17_Cmult29} {iopath_Amult17_Cmult30} {iopath_Amult17_Cmult31} {iopath_Amult17_Cmult32} {iopath_Amult17_Cmult33} {iopath_Amult17_Cmult34} {iopath_Amult17_Cmult35} {iopath_Amult17_Cmult36} {iopath_Amult17_Cmult37} {iopath_Amult17_Cmult38} {iopath_Amult17_Cmult39} {iopath_Amult17_Cmult40} {iopath_Amult17_Cmult41} {iopath_Amult17_Cmult42} {iopath_Amult17_Cmult43} {iopath_Amult17_Cmult44} {iopath_Amult17_Cmult45} {iopath_Amult17_Cmult46} {iopath_Amult17_Cmult47} {iopath_Amult17_Cmult48} {iopath_Amult17_Cmult49} {iopath_Amult17_Cmult50} {iopath_Amult17_Cmult51} {iopath_Amult17_Cmult52} {iopath_Amult17_Cmult53} {iopath_Amult17_Cmult54} {iopath_Amult17_Cmult55} {iopath_Amult17_Cmult56} {iopath_Amult17_Cmult57} {iopath_Amult17_Cmult58} {iopath_Amult17_Cmult59} {iopath_Amult17_Cmult60} {iopath_Amult17_Cmult61} {iopath_Amult17_Cmult62} {iopath_Amult17_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult18_Cmult18} {iopath_Amult18_Cmult19} {iopath_Amult18_Cmult20} {iopath_Amult18_Cmult21} {iopath_Amult18_Cmult22} {iopath_Amult18_Cmult23} {iopath_Amult18_Cmult24} {iopath_Amult18_Cmult25} {iopath_Amult18_Cmult26} {iopath_Amult18_Cmult27} {iopath_Amult18_Cmult28} {iopath_Amult18_Cmult29} {iopath_Amult18_Cmult30} {iopath_Amult18_Cmult31} {iopath_Amult18_Cmult32} {iopath_Amult18_Cmult33} {iopath_Amult18_Cmult34} {iopath_Amult18_Cmult35} {iopath_Amult18_Cmult36} {iopath_Amult18_Cmult37} {iopath_Amult18_Cmult38} {iopath_Amult18_Cmult39} {iopath_Amult18_Cmult40} {iopath_Amult18_Cmult41} {iopath_Amult18_Cmult42} {iopath_Amult18_Cmult43} {iopath_Amult18_Cmult44} {iopath_Amult18_Cmult45} {iopath_Amult18_Cmult46} {iopath_Amult18_Cmult47} {iopath_Amult18_Cmult48} {iopath_Amult18_Cmult49} {iopath_Amult18_Cmult50} {iopath_Amult18_Cmult51} {iopath_Amult18_Cmult52} {iopath_Amult18_Cmult53} {iopath_Amult18_Cmult54} {iopath_Amult18_Cmult55} {iopath_Amult18_Cmult56} {iopath_Amult18_Cmult57} {iopath_Amult18_Cmult58} {iopath_Amult18_Cmult59} {iopath_Amult18_Cmult60} {iopath_Amult18_Cmult61} {iopath_Amult18_Cmult62} {iopath_Amult18_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult19_Cmult19} {iopath_Amult19_Cmult20} {iopath_Amult19_Cmult21} {iopath_Amult19_Cmult22} {iopath_Amult19_Cmult23} {iopath_Amult19_Cmult24} {iopath_Amult19_Cmult25} {iopath_Amult19_Cmult26} {iopath_Amult19_Cmult27} {iopath_Amult19_Cmult28} {iopath_Amult19_Cmult29} {iopath_Amult19_Cmult30} {iopath_Amult19_Cmult31} {iopath_Amult19_Cmult32} {iopath_Amult19_Cmult33} {iopath_Amult19_Cmult34} {iopath_Amult19_Cmult35} {iopath_Amult19_Cmult36} {iopath_Amult19_Cmult37} {iopath_Amult19_Cmult38} {iopath_Amult19_Cmult39} {iopath_Amult19_Cmult40} {iopath_Amult19_Cmult41} {iopath_Amult19_Cmult42} {iopath_Amult19_Cmult43} {iopath_Amult19_Cmult44} {iopath_Amult19_Cmult45} {iopath_Amult19_Cmult46} {iopath_Amult19_Cmult47} {iopath_Amult19_Cmult48} {iopath_Amult19_Cmult49} {iopath_Amult19_Cmult50} {iopath_Amult19_Cmult51} {iopath_Amult19_Cmult52} {iopath_Amult19_Cmult53} {iopath_Amult19_Cmult54} {iopath_Amult19_Cmult55} {iopath_Amult19_Cmult56} {iopath_Amult19_Cmult57} {iopath_Amult19_Cmult58} {iopath_Amult19_Cmult59} {iopath_Amult19_Cmult60} {iopath_Amult19_Cmult61} {iopath_Amult19_Cmult62} {iopath_Amult19_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult20_Cmult20} {iopath_Amult20_Cmult21} {iopath_Amult20_Cmult22} {iopath_Amult20_Cmult23} {iopath_Amult20_Cmult24} {iopath_Amult20_Cmult25} {iopath_Amult20_Cmult26} {iopath_Amult20_Cmult27} {iopath_Amult20_Cmult28} {iopath_Amult20_Cmult29} {iopath_Amult20_Cmult30} {iopath_Amult20_Cmult31} {iopath_Amult20_Cmult32} {iopath_Amult20_Cmult33} {iopath_Amult20_Cmult34} {iopath_Amult20_Cmult35} {iopath_Amult20_Cmult36} {iopath_Amult20_Cmult37} {iopath_Amult20_Cmult38} {iopath_Amult20_Cmult39} {iopath_Amult20_Cmult40} {iopath_Amult20_Cmult41} {iopath_Amult20_Cmult42} {iopath_Amult20_Cmult43} {iopath_Amult20_Cmult44} {iopath_Amult20_Cmult45} {iopath_Amult20_Cmult46} {iopath_Amult20_Cmult47} {iopath_Amult20_Cmult48} {iopath_Amult20_Cmult49} {iopath_Amult20_Cmult50} {iopath_Amult20_Cmult51} {iopath_Amult20_Cmult52} {iopath_Amult20_Cmult53} {iopath_Amult20_Cmult54} {iopath_Amult20_Cmult55} {iopath_Amult20_Cmult56} {iopath_Amult20_Cmult57} {iopath_Amult20_Cmult58} {iopath_Amult20_Cmult59} {iopath_Amult20_Cmult60} {iopath_Amult20_Cmult61} {iopath_Amult20_Cmult62} {iopath_Amult20_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult21_Cmult21} {iopath_Amult21_Cmult22} {iopath_Amult21_Cmult23} {iopath_Amult21_Cmult24} {iopath_Amult21_Cmult25} {iopath_Amult21_Cmult26} {iopath_Amult21_Cmult27} {iopath_Amult21_Cmult28} {iopath_Amult21_Cmult29} {iopath_Amult21_Cmult30} {iopath_Amult21_Cmult31} {iopath_Amult21_Cmult32} {iopath_Amult21_Cmult33} {iopath_Amult21_Cmult34} {iopath_Amult21_Cmult35} {iopath_Amult21_Cmult36} {iopath_Amult21_Cmult37} {iopath_Amult21_Cmult38} {iopath_Amult21_Cmult39} {iopath_Amult21_Cmult40} {iopath_Amult21_Cmult41} {iopath_Amult21_Cmult42} {iopath_Amult21_Cmult43} {iopath_Amult21_Cmult44} {iopath_Amult21_Cmult45} {iopath_Amult21_Cmult46} {iopath_Amult21_Cmult47} {iopath_Amult21_Cmult48} {iopath_Amult21_Cmult49} {iopath_Amult21_Cmult50} {iopath_Amult21_Cmult51} {iopath_Amult21_Cmult52} {iopath_Amult21_Cmult53} {iopath_Amult21_Cmult54} {iopath_Amult21_Cmult55} {iopath_Amult21_Cmult56} {iopath_Amult21_Cmult57} {iopath_Amult21_Cmult58} {iopath_Amult21_Cmult59} {iopath_Amult21_Cmult60} {iopath_Amult21_Cmult61} {iopath_Amult21_Cmult62} {iopath_Amult21_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult22_Cmult22} {iopath_Amult22_Cmult23} {iopath_Amult22_Cmult24} {iopath_Amult22_Cmult25} {iopath_Amult22_Cmult26} {iopath_Amult22_Cmult27} {iopath_Amult22_Cmult28} {iopath_Amult22_Cmult29} {iopath_Amult22_Cmult30} {iopath_Amult22_Cmult31} {iopath_Amult22_Cmult32} {iopath_Amult22_Cmult33} {iopath_Amult22_Cmult34} {iopath_Amult22_Cmult35} {iopath_Amult22_Cmult36} {iopath_Amult22_Cmult37} {iopath_Amult22_Cmult38} {iopath_Amult22_Cmult39} {iopath_Amult22_Cmult40} {iopath_Amult22_Cmult41} {iopath_Amult22_Cmult42} {iopath_Amult22_Cmult43} {iopath_Amult22_Cmult44} {iopath_Amult22_Cmult45} {iopath_Amult22_Cmult46} {iopath_Amult22_Cmult47} {iopath_Amult22_Cmult48} {iopath_Amult22_Cmult49} {iopath_Amult22_Cmult50} {iopath_Amult22_Cmult51} {iopath_Amult22_Cmult52} {iopath_Amult22_Cmult53} {iopath_Amult22_Cmult54} {iopath_Amult22_Cmult55} {iopath_Amult22_Cmult56} {iopath_Amult22_Cmult57} {iopath_Amult22_Cmult58} {iopath_Amult22_Cmult59} {iopath_Amult22_Cmult60} {iopath_Amult22_Cmult61} {iopath_Amult22_Cmult62} {iopath_Amult22_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult23_Cmult23} {iopath_Amult23_Cmult24} {iopath_Amult23_Cmult25} {iopath_Amult23_Cmult26} {iopath_Amult23_Cmult27} {iopath_Amult23_Cmult28} {iopath_Amult23_Cmult29} {iopath_Amult23_Cmult30} {iopath_Amult23_Cmult31} {iopath_Amult23_Cmult32} {iopath_Amult23_Cmult33} {iopath_Amult23_Cmult34} {iopath_Amult23_Cmult35} {iopath_Amult23_Cmult36} {iopath_Amult23_Cmult37} {iopath_Amult23_Cmult38} {iopath_Amult23_Cmult39} {iopath_Amult23_Cmult40} {iopath_Amult23_Cmult41} {iopath_Amult23_Cmult42} {iopath_Amult23_Cmult43} {iopath_Amult23_Cmult44} {iopath_Amult23_Cmult45} {iopath_Amult23_Cmult46} {iopath_Amult23_Cmult47} {iopath_Amult23_Cmult48} {iopath_Amult23_Cmult49} {iopath_Amult23_Cmult50} {iopath_Amult23_Cmult51} {iopath_Amult23_Cmult52} {iopath_Amult23_Cmult53} {iopath_Amult23_Cmult54} {iopath_Amult23_Cmult55} {iopath_Amult23_Cmult56} {iopath_Amult23_Cmult57} {iopath_Amult23_Cmult58} {iopath_Amult23_Cmult59} {iopath_Amult23_Cmult60} {iopath_Amult23_Cmult61} {iopath_Amult23_Cmult62} {iopath_Amult23_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult24_Cmult24} {iopath_Amult24_Cmult25} {iopath_Amult24_Cmult26} {iopath_Amult24_Cmult27} {iopath_Amult24_Cmult28} {iopath_Amult24_Cmult29} {iopath_Amult24_Cmult30} {iopath_Amult24_Cmult31} {iopath_Amult24_Cmult32} {iopath_Amult24_Cmult33} {iopath_Amult24_Cmult34} {iopath_Amult24_Cmult35} {iopath_Amult24_Cmult36} {iopath_Amult24_Cmult37} {iopath_Amult24_Cmult38} {iopath_Amult24_Cmult39} {iopath_Amult24_Cmult40} {iopath_Amult24_Cmult41} {iopath_Amult24_Cmult42} {iopath_Amult24_Cmult43} {iopath_Amult24_Cmult44} {iopath_Amult24_Cmult45} {iopath_Amult24_Cmult46} {iopath_Amult24_Cmult47} {iopath_Amult24_Cmult48} {iopath_Amult24_Cmult49} {iopath_Amult24_Cmult50} {iopath_Amult24_Cmult51} {iopath_Amult24_Cmult52} {iopath_Amult24_Cmult53} {iopath_Amult24_Cmult54} {iopath_Amult24_Cmult55} {iopath_Amult24_Cmult56} {iopath_Amult24_Cmult57} {iopath_Amult24_Cmult58} {iopath_Amult24_Cmult59} {iopath_Amult24_Cmult60} {iopath_Amult24_Cmult61} {iopath_Amult24_Cmult62} {iopath_Amult24_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult25_Cmult25} {iopath_Amult25_Cmult26} {iopath_Amult25_Cmult27} {iopath_Amult25_Cmult28} {iopath_Amult25_Cmult29} {iopath_Amult25_Cmult30} {iopath_Amult25_Cmult31} {iopath_Amult25_Cmult32} {iopath_Amult25_Cmult33} {iopath_Amult25_Cmult34} {iopath_Amult25_Cmult35} {iopath_Amult25_Cmult36} {iopath_Amult25_Cmult37} {iopath_Amult25_Cmult38} {iopath_Amult25_Cmult39} {iopath_Amult25_Cmult40} {iopath_Amult25_Cmult41} {iopath_Amult25_Cmult42} {iopath_Amult25_Cmult43} {iopath_Amult25_Cmult44} {iopath_Amult25_Cmult45} {iopath_Amult25_Cmult46} {iopath_Amult25_Cmult47} {iopath_Amult25_Cmult48} {iopath_Amult25_Cmult49} {iopath_Amult25_Cmult50} {iopath_Amult25_Cmult51} {iopath_Amult25_Cmult52} {iopath_Amult25_Cmult53} {iopath_Amult25_Cmult54} {iopath_Amult25_Cmult55} {iopath_Amult25_Cmult56} {iopath_Amult25_Cmult57} {iopath_Amult25_Cmult58} {iopath_Amult25_Cmult59} {iopath_Amult25_Cmult60} {iopath_Amult25_Cmult61} {iopath_Amult25_Cmult62} {iopath_Amult25_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult26_Cmult26} {iopath_Amult26_Cmult27} {iopath_Amult26_Cmult28} {iopath_Amult26_Cmult29} {iopath_Amult26_Cmult30} {iopath_Amult26_Cmult31} {iopath_Amult26_Cmult32} {iopath_Amult26_Cmult33} {iopath_Amult26_Cmult34} {iopath_Amult26_Cmult35} {iopath_Amult26_Cmult36} {iopath_Amult26_Cmult37} {iopath_Amult26_Cmult38} {iopath_Amult26_Cmult39} {iopath_Amult26_Cmult40} {iopath_Amult26_Cmult41} {iopath_Amult26_Cmult42} {iopath_Amult26_Cmult43} {iopath_Amult26_Cmult44} {iopath_Amult26_Cmult45} {iopath_Amult26_Cmult46} {iopath_Amult26_Cmult47} {iopath_Amult26_Cmult48} {iopath_Amult26_Cmult49} {iopath_Amult26_Cmult50} {iopath_Amult26_Cmult51} {iopath_Amult26_Cmult52} {iopath_Amult26_Cmult53} {iopath_Amult26_Cmult54} {iopath_Amult26_Cmult55} {iopath_Amult26_Cmult56} {iopath_Amult26_Cmult57} {iopath_Amult26_Cmult58} {iopath_Amult26_Cmult59} {iopath_Amult26_Cmult60} {iopath_Amult26_Cmult61} {iopath_Amult26_Cmult62} {iopath_Amult26_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult27_Cmult27} {iopath_Amult27_Cmult28} {iopath_Amult27_Cmult29} {iopath_Amult27_Cmult30} {iopath_Amult27_Cmult31} {iopath_Amult27_Cmult32} {iopath_Amult27_Cmult33} {iopath_Amult27_Cmult34} {iopath_Amult27_Cmult35} {iopath_Amult27_Cmult36} {iopath_Amult27_Cmult37} {iopath_Amult27_Cmult38} {iopath_Amult27_Cmult39} {iopath_Amult27_Cmult40} {iopath_Amult27_Cmult41} {iopath_Amult27_Cmult42} {iopath_Amult27_Cmult43} {iopath_Amult27_Cmult44} {iopath_Amult27_Cmult45} {iopath_Amult27_Cmult46} {iopath_Amult27_Cmult47} {iopath_Amult27_Cmult48} {iopath_Amult27_Cmult49} {iopath_Amult27_Cmult50} {iopath_Amult27_Cmult51} {iopath_Amult27_Cmult52} {iopath_Amult27_Cmult53} {iopath_Amult27_Cmult54} {iopath_Amult27_Cmult55} {iopath_Amult27_Cmult56} {iopath_Amult27_Cmult57} {iopath_Amult27_Cmult58} {iopath_Amult27_Cmult59} {iopath_Amult27_Cmult60} {iopath_Amult27_Cmult61} {iopath_Amult27_Cmult62} {iopath_Amult27_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult28_Cmult28} {iopath_Amult28_Cmult29} {iopath_Amult28_Cmult30} {iopath_Amult28_Cmult31} {iopath_Amult28_Cmult32} {iopath_Amult28_Cmult33} {iopath_Amult28_Cmult34} {iopath_Amult28_Cmult35} {iopath_Amult28_Cmult36} {iopath_Amult28_Cmult37} {iopath_Amult28_Cmult38} {iopath_Amult28_Cmult39} {iopath_Amult28_Cmult40} {iopath_Amult28_Cmult41} {iopath_Amult28_Cmult42} {iopath_Amult28_Cmult43} {iopath_Amult28_Cmult44} {iopath_Amult28_Cmult45} {iopath_Amult28_Cmult46} {iopath_Amult28_Cmult47} {iopath_Amult28_Cmult48} {iopath_Amult28_Cmult49} {iopath_Amult28_Cmult50} {iopath_Amult28_Cmult51} {iopath_Amult28_Cmult52} {iopath_Amult28_Cmult53} {iopath_Amult28_Cmult54} {iopath_Amult28_Cmult55} {iopath_Amult28_Cmult56} {iopath_Amult28_Cmult57} {iopath_Amult28_Cmult58} {iopath_Amult28_Cmult59} {iopath_Amult28_Cmult60} {iopath_Amult28_Cmult61} {iopath_Amult28_Cmult62} {iopath_Amult28_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult29_Cmult29} {iopath_Amult29_Cmult30} {iopath_Amult29_Cmult31} {iopath_Amult29_Cmult32} {iopath_Amult29_Cmult33} {iopath_Amult29_Cmult34} {iopath_Amult29_Cmult35} {iopath_Amult29_Cmult36} {iopath_Amult29_Cmult37} {iopath_Amult29_Cmult38} {iopath_Amult29_Cmult39} {iopath_Amult29_Cmult40} {iopath_Amult29_Cmult41} {iopath_Amult29_Cmult42} {iopath_Amult29_Cmult43} {iopath_Amult29_Cmult44} {iopath_Amult29_Cmult45} {iopath_Amult29_Cmult46} {iopath_Amult29_Cmult47} {iopath_Amult29_Cmult48} {iopath_Amult29_Cmult49} {iopath_Amult29_Cmult50} {iopath_Amult29_Cmult51} {iopath_Amult29_Cmult52} {iopath_Amult29_Cmult53} {iopath_Amult29_Cmult54} {iopath_Amult29_Cmult55} {iopath_Amult29_Cmult56} {iopath_Amult29_Cmult57} {iopath_Amult29_Cmult58} {iopath_Amult29_Cmult59} {iopath_Amult29_Cmult60} {iopath_Amult29_Cmult61} {iopath_Amult29_Cmult62} {iopath_Amult29_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult30_Cmult30} {iopath_Amult30_Cmult31} {iopath_Amult30_Cmult32} {iopath_Amult30_Cmult33} {iopath_Amult30_Cmult34} {iopath_Amult30_Cmult35} {iopath_Amult30_Cmult36} {iopath_Amult30_Cmult37} {iopath_Amult30_Cmult38} {iopath_Amult30_Cmult39} {iopath_Amult30_Cmult40} {iopath_Amult30_Cmult41} {iopath_Amult30_Cmult42} {iopath_Amult30_Cmult43} {iopath_Amult30_Cmult44} {iopath_Amult30_Cmult45} {iopath_Amult30_Cmult46} {iopath_Amult30_Cmult47} {iopath_Amult30_Cmult48} {iopath_Amult30_Cmult49} {iopath_Amult30_Cmult50} {iopath_Amult30_Cmult51} {iopath_Amult30_Cmult52} {iopath_Amult30_Cmult53} {iopath_Amult30_Cmult54} {iopath_Amult30_Cmult55} {iopath_Amult30_Cmult56} {iopath_Amult30_Cmult57} {iopath_Amult30_Cmult58} {iopath_Amult30_Cmult59} {iopath_Amult30_Cmult60} {iopath_Amult30_Cmult61} {iopath_Amult30_Cmult62} {iopath_Amult30_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult31_Cmult31} {iopath_Amult31_Cmult32} {iopath_Amult31_Cmult33} {iopath_Amult31_Cmult34} {iopath_Amult31_Cmult35} {iopath_Amult31_Cmult36} {iopath_Amult31_Cmult37} {iopath_Amult31_Cmult38} {iopath_Amult31_Cmult39} {iopath_Amult31_Cmult40} {iopath_Amult31_Cmult41} {iopath_Amult31_Cmult42} {iopath_Amult31_Cmult43} {iopath_Amult31_Cmult44} {iopath_Amult31_Cmult45} {iopath_Amult31_Cmult46} {iopath_Amult31_Cmult47} {iopath_Amult31_Cmult48} {iopath_Amult31_Cmult49} {iopath_Amult31_Cmult50} {iopath_Amult31_Cmult51} {iopath_Amult31_Cmult52} {iopath_Amult31_Cmult53} {iopath_Amult31_Cmult54} {iopath_Amult31_Cmult55} {iopath_Amult31_Cmult56} {iopath_Amult31_Cmult57} {iopath_Amult31_Cmult58} {iopath_Amult31_Cmult59} {iopath_Amult31_Cmult60} {iopath_Amult31_Cmult61} {iopath_Amult31_Cmult62} {iopath_Amult31_Cmult63} "*)
	(* DELAY_MATRIX_Valid_mult="1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 "*)
	(* DELAY_MATRIX_sel_mul_32x32="1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 "*)
	output reg  [63:0] Cmult;
	input wire         sel_mul_32x32;

`ifdef GSIM
    specify
		(Amult[0]  => Cmult[0]) = "";
		(Amult[1]  => Cmult[0]) = "";
		(Amult[2]  => Cmult[0]) = "";
		(Amult[3]  => Cmult[0]) = "";
		(Amult[4]  => Cmult[0]) = "";
		(Amult[5]  => Cmult[0]) = "";
		(Amult[6]  => Cmult[0]) = "";
		(Amult[7]  => Cmult[0]) = "";
		(Amult[8]  => Cmult[0]) = "";
		(Amult[9]  => Cmult[0]) = "";
		(Amult[10] => Cmult[0]) = "";
		(Amult[11] => Cmult[0]) = "";
		(Amult[12] => Cmult[0]) = "";
		(Amult[13] => Cmult[0]) = "";
		(Amult[14] => Cmult[0]) = "";
		(Amult[15] => Cmult[0]) = "";
		(Amult[16] => Cmult[0]) = "";
		(Amult[17] => Cmult[0]) = "";
		(Amult[18] => Cmult[0]) = "";
		(Amult[19] => Cmult[0]) = "";
		(Amult[20] => Cmult[0]) = "";
		(Amult[21] => Cmult[0]) = "";
		(Amult[22] => Cmult[0]) = "";
		(Amult[23] => Cmult[0]) = "";
		(Amult[24] => Cmult[0]) = "";
		(Amult[25] => Cmult[0]) = "";
		(Amult[26] => Cmult[0]) = "";
		(Amult[27] => Cmult[0]) = "";
		(Amult[28] => Cmult[0]) = "";
		(Amult[29] => Cmult[0]) = "";
		(Amult[30] => Cmult[0]) = "";
		(Amult[31] => Cmult[0]) = "";
		(Bmult[0]  => Cmult[0]) = "";
		(Bmult[1]  => Cmult[0]) = "";
		(Bmult[2]  => Cmult[0]) = "";
		(Bmult[3]  => Cmult[0]) = "";
		(Bmult[4]  => Cmult[0]) = "";
		(Bmult[5]  => Cmult[0]) = "";
		(Bmult[6]  => Cmult[0]) = "";
		(Bmult[7]  => Cmult[0]) = "";
		(Bmult[8]  => Cmult[0]) = "";
		(Bmult[9]  => Cmult[0]) = "";
		(Bmult[10] => Cmult[0]) = "";
		(Bmult[11] => Cmult[0]) = "";
		(Bmult[12] => Cmult[0]) = "";
		(Bmult[13] => Cmult[0]) = "";
		(Bmult[14] => Cmult[0]) = "";
		(Bmult[15] => Cmult[0]) = "";
		(Bmult[16] => Cmult[0]) = "";
		(Bmult[17] => Cmult[0]) = "";
		(Bmult[18] => Cmult[0]) = "";
		(Bmult[19] => Cmult[0]) = "";
		(Bmult[20] => Cmult[0]) = "";
		(Bmult[21] => Cmult[0]) = "";
		(Bmult[22] => Cmult[0]) = "";
		(Bmult[23] => Cmult[0]) = "";
		(Bmult[24] => Cmult[0]) = "";
		(Bmult[25] => Cmult[0]) = "";
		(Bmult[26] => Cmult[0]) = "";
		(Bmult[27] => Cmult[0]) = "";
		(Bmult[28] => Cmult[0]) = "";
		(Bmult[29] => Cmult[0]) = "";
		(Bmult[30] => Cmult[0]) = "";
		(Bmult[31] => Cmult[0]) = "";		
		(Valid_mult[0] => Cmult[0]) = "";
		(Valid_mult[1] => Cmult[0]) = "";
		(sel_mul_32x32 => Cmult[0]) = "";
		(Amult[0]  => Cmult[1]) = "";
		(Amult[1]  => Cmult[1]) = "";
		(Amult[2]  => Cmult[1]) = "";
		(Amult[3]  => Cmult[1]) = "";
		(Amult[4]  => Cmult[1]) = "";
		(Amult[5]  => Cmult[1]) = "";
		(Amult[6]  => Cmult[1]) = "";
		(Amult[7]  => Cmult[1]) = "";
		(Amult[8]  => Cmult[1]) = "";
		(Amult[9]  => Cmult[1]) = "";
		(Amult[10] => Cmult[1]) = "";
		(Amult[11] => Cmult[1]) = "";
		(Amult[12] => Cmult[1]) = "";
		(Amult[13] => Cmult[1]) = "";
		(Amult[14] => Cmult[1]) = "";
		(Amult[15] => Cmult[1]) = "";
		(Amult[16] => Cmult[1]) = "";
		(Amult[17] => Cmult[1]) = "";
		(Amult[18] => Cmult[1]) = "";
		(Amult[19] => Cmult[1]) = "";
		(Amult[20] => Cmult[1]) = "";
		(Amult[21] => Cmult[1]) = "";
		(Amult[22] => Cmult[1]) = "";
		(Amult[23] => Cmult[1]) = "";
		(Amult[24] => Cmult[1]) = "";
		(Amult[25] => Cmult[1]) = "";
		(Amult[26] => Cmult[1]) = "";
		(Amult[27] => Cmult[1]) = "";
		(Amult[28] => Cmult[1]) = "";
		(Amult[29] => Cmult[1]) = "";
		(Amult[30] => Cmult[1]) = "";
		(Amult[31] => Cmult[1]) = "";
		(Bmult[0]  => Cmult[1]) = "";
		(Bmult[1]  => Cmult[1]) = "";
		(Bmult[2]  => Cmult[1]) = "";
		(Bmult[3]  => Cmult[1]) = "";
		(Bmult[4]  => Cmult[1]) = "";
		(Bmult[5]  => Cmult[1]) = "";
		(Bmult[6]  => Cmult[1]) = "";
		(Bmult[7]  => Cmult[1]) = "";
		(Bmult[8]  => Cmult[1]) = "";
		(Bmult[9]  => Cmult[1]) = "";
		(Bmult[10] => Cmult[1]) = "";
		(Bmult[11] => Cmult[1]) = "";
		(Bmult[12] => Cmult[1]) = "";
		(Bmult[13] => Cmult[1]) = "";
		(Bmult[14] => Cmult[1]) = "";
		(Bmult[15] => Cmult[1]) = "";
		(Bmult[16] => Cmult[1]) = "";
		(Bmult[17] => Cmult[1]) = "";
		(Bmult[18] => Cmult[1]) = "";
		(Bmult[19] => Cmult[1]) = "";
		(Bmult[20] => Cmult[1]) = "";
		(Bmult[21] => Cmult[1]) = "";
		(Bmult[22] => Cmult[1]) = "";
		(Bmult[23] => Cmult[1]) = "";
		(Bmult[24] => Cmult[1]) = "";
		(Bmult[25] => Cmult[1]) = "";
		(Bmult[26] => Cmult[1]) = "";
		(Bmult[27] => Cmult[1]) = "";
		(Bmult[28] => Cmult[1]) = "";
		(Bmult[29] => Cmult[1]) = "";
		(Bmult[30] => Cmult[1]) = "";
		(Bmult[31] => Cmult[1]) = "";		
		(Valid_mult[0] => Cmult[1]) = "";
		(Valid_mult[1] => Cmult[1]) = "";
		(sel_mul_32x32 => Cmult[1]) = "";
		(Amult[0]  => Cmult[2]) = "";
		(Amult[1]  => Cmult[2]) = "";
		(Amult[2]  => Cmult[2]) = "";
		(Amult[3]  => Cmult[2]) = "";
		(Amult[4]  => Cmult[2]) = "";
		(Amult[5]  => Cmult[2]) = "";
		(Amult[6]  => Cmult[2]) = "";
		(Amult[7]  => Cmult[2]) = "";
		(Amult[8]  => Cmult[2]) = "";
		(Amult[9]  => Cmult[2]) = "";
		(Amult[10] => Cmult[2]) = "";
		(Amult[11] => Cmult[2]) = "";
		(Amult[12] => Cmult[2]) = "";
		(Amult[13] => Cmult[2]) = "";
		(Amult[14] => Cmult[2]) = "";
		(Amult[15] => Cmult[2]) = "";
		(Amult[16] => Cmult[2]) = "";
		(Amult[17] => Cmult[2]) = "";
		(Amult[18] => Cmult[2]) = "";
		(Amult[19] => Cmult[2]) = "";
		(Amult[20] => Cmult[2]) = "";
		(Amult[21] => Cmult[2]) = "";
		(Amult[22] => Cmult[2]) = "";
		(Amult[23] => Cmult[2]) = "";
		(Amult[24] => Cmult[2]) = "";
		(Amult[25] => Cmult[2]) = "";
		(Amult[26] => Cmult[2]) = "";
		(Amult[27] => Cmult[2]) = "";
		(Amult[28] => Cmult[2]) = "";
		(Amult[29] => Cmult[2]) = "";
		(Amult[30] => Cmult[2]) = "";
		(Amult[31] => Cmult[2]) = "";
		(Bmult[0]  => Cmult[2]) = "";
		(Bmult[1]  => Cmult[2]) = "";
		(Bmult[2]  => Cmult[2]) = "";
		(Bmult[3]  => Cmult[2]) = "";
		(Bmult[4]  => Cmult[2]) = "";
		(Bmult[5]  => Cmult[2]) = "";
		(Bmult[6]  => Cmult[2]) = "";
		(Bmult[7]  => Cmult[2]) = "";
		(Bmult[8]  => Cmult[2]) = "";
		(Bmult[9]  => Cmult[2]) = "";
		(Bmult[10] => Cmult[2]) = "";
		(Bmult[11] => Cmult[2]) = "";
		(Bmult[12] => Cmult[2]) = "";
		(Bmult[13] => Cmult[2]) = "";
		(Bmult[14] => Cmult[2]) = "";
		(Bmult[15] => Cmult[2]) = "";
		(Bmult[16] => Cmult[2]) = "";
		(Bmult[17] => Cmult[2]) = "";
		(Bmult[18] => Cmult[2]) = "";
		(Bmult[19] => Cmult[2]) = "";
		(Bmult[20] => Cmult[2]) = "";
		(Bmult[21] => Cmult[2]) = "";
		(Bmult[22] => Cmult[2]) = "";
		(Bmult[23] => Cmult[2]) = "";
		(Bmult[24] => Cmult[2]) = "";
		(Bmult[25] => Cmult[2]) = "";
		(Bmult[26] => Cmult[2]) = "";
		(Bmult[27] => Cmult[2]) = "";
		(Bmult[28] => Cmult[2]) = "";
		(Bmult[29] => Cmult[2]) = "";
		(Bmult[30] => Cmult[2]) = "";
		(Bmult[31] => Cmult[2]) = "";		
		(Valid_mult[0] => Cmult[2]) = "";
		(Valid_mult[1] => Cmult[2]) = "";
		(sel_mul_32x32 => Cmult[2]) = "";
		(Amult[0]  => Cmult[3]) = "";
		(Amult[1]  => Cmult[3]) = "";
		(Amult[2]  => Cmult[3]) = "";
		(Amult[3]  => Cmult[3]) = "";
		(Amult[4]  => Cmult[3]) = "";
		(Amult[5]  => Cmult[3]) = "";
		(Amult[6]  => Cmult[3]) = "";
		(Amult[7]  => Cmult[3]) = "";
		(Amult[8]  => Cmult[3]) = "";
		(Amult[9]  => Cmult[3]) = "";
		(Amult[10] => Cmult[3]) = "";
		(Amult[11] => Cmult[3]) = "";
		(Amult[12] => Cmult[3]) = "";
		(Amult[13] => Cmult[3]) = "";
		(Amult[14] => Cmult[3]) = "";
		(Amult[15] => Cmult[3]) = "";
		(Amult[16] => Cmult[3]) = "";
		(Amult[17] => Cmult[3]) = "";
		(Amult[18] => Cmult[3]) = "";
		(Amult[19] => Cmult[3]) = "";
		(Amult[20] => Cmult[3]) = "";
		(Amult[21] => Cmult[3]) = "";
		(Amult[22] => Cmult[3]) = "";
		(Amult[23] => Cmult[3]) = "";
		(Amult[24] => Cmult[3]) = "";
		(Amult[25] => Cmult[3]) = "";
		(Amult[26] => Cmult[3]) = "";
		(Amult[27] => Cmult[3]) = "";
		(Amult[28] => Cmult[3]) = "";
		(Amult[29] => Cmult[3]) = "";
		(Amult[30] => Cmult[3]) = "";
		(Amult[31] => Cmult[3]) = "";
		(Bmult[0]  => Cmult[3]) = "";
		(Bmult[1]  => Cmult[3]) = "";
		(Bmult[2]  => Cmult[3]) = "";
		(Bmult[3]  => Cmult[3]) = "";
		(Bmult[4]  => Cmult[3]) = "";
		(Bmult[5]  => Cmult[3]) = "";
		(Bmult[6]  => Cmult[3]) = "";
		(Bmult[7]  => Cmult[3]) = "";
		(Bmult[8]  => Cmult[3]) = "";
		(Bmult[9]  => Cmult[3]) = "";
		(Bmult[10] => Cmult[3]) = "";
		(Bmult[11] => Cmult[3]) = "";
		(Bmult[12] => Cmult[3]) = "";
		(Bmult[13] => Cmult[3]) = "";
		(Bmult[14] => Cmult[3]) = "";
		(Bmult[15] => Cmult[3]) = "";
		(Bmult[16] => Cmult[3]) = "";
		(Bmult[17] => Cmult[3]) = "";
		(Bmult[18] => Cmult[3]) = "";
		(Bmult[19] => Cmult[3]) = "";
		(Bmult[20] => Cmult[3]) = "";
		(Bmult[21] => Cmult[3]) = "";
		(Bmult[22] => Cmult[3]) = "";
		(Bmult[23] => Cmult[3]) = "";
		(Bmult[24] => Cmult[3]) = "";
		(Bmult[25] => Cmult[3]) = "";
		(Bmult[26] => Cmult[3]) = "";
		(Bmult[27] => Cmult[3]) = "";
		(Bmult[28] => Cmult[3]) = "";
		(Bmult[29] => Cmult[3]) = "";
		(Bmult[30] => Cmult[3]) = "";
		(Bmult[31] => Cmult[3]) = "";		
		(Valid_mult[0] => Cmult[3]) = "";
		(Valid_mult[1] => Cmult[3]) = "";
		(sel_mul_32x32 => Cmult[3]) = "";
		(Amult[0]  => Cmult[4]) = "";
		(Amult[1]  => Cmult[4]) = "";
		(Amult[2]  => Cmult[4]) = "";
		(Amult[3]  => Cmult[4]) = "";
		(Amult[4]  => Cmult[4]) = "";
		(Amult[5]  => Cmult[4]) = "";
		(Amult[6]  => Cmult[4]) = "";
		(Amult[7]  => Cmult[4]) = "";
		(Amult[8]  => Cmult[4]) = "";
		(Amult[9]  => Cmult[4]) = "";
		(Amult[10] => Cmult[4]) = "";
		(Amult[11] => Cmult[4]) = "";
		(Amult[12] => Cmult[4]) = "";
		(Amult[13] => Cmult[4]) = "";
		(Amult[14] => Cmult[4]) = "";
		(Amult[15] => Cmult[4]) = "";
		(Amult[16] => Cmult[4]) = "";
		(Amult[17] => Cmult[4]) = "";
		(Amult[18] => Cmult[4]) = "";
		(Amult[19] => Cmult[4]) = "";
		(Amult[20] => Cmult[4]) = "";
		(Amult[21] => Cmult[4]) = "";
		(Amult[22] => Cmult[4]) = "";
		(Amult[23] => Cmult[4]) = "";
		(Amult[24] => Cmult[4]) = "";
		(Amult[25] => Cmult[4]) = "";
		(Amult[26] => Cmult[4]) = "";
		(Amult[27] => Cmult[4]) = "";
		(Amult[28] => Cmult[4]) = "";
		(Amult[29] => Cmult[4]) = "";
		(Amult[30] => Cmult[4]) = "";
		(Amult[31] => Cmult[4]) = "";
		(Bmult[0]  => Cmult[4]) = "";
		(Bmult[1]  => Cmult[4]) = "";
		(Bmult[2]  => Cmult[4]) = "";
		(Bmult[3]  => Cmult[4]) = "";
		(Bmult[4]  => Cmult[4]) = "";
		(Bmult[5]  => Cmult[4]) = "";
		(Bmult[6]  => Cmult[4]) = "";
		(Bmult[7]  => Cmult[4]) = "";
		(Bmult[8]  => Cmult[4]) = "";
		(Bmult[9]  => Cmult[4]) = "";
		(Bmult[10] => Cmult[4]) = "";
		(Bmult[11] => Cmult[4]) = "";
		(Bmult[12] => Cmult[4]) = "";
		(Bmult[13] => Cmult[4]) = "";
		(Bmult[14] => Cmult[4]) = "";
		(Bmult[15] => Cmult[4]) = "";
		(Bmult[16] => Cmult[4]) = "";
		(Bmult[17] => Cmult[4]) = "";
		(Bmult[18] => Cmult[4]) = "";
		(Bmult[19] => Cmult[4]) = "";
		(Bmult[20] => Cmult[4]) = "";
		(Bmult[21] => Cmult[4]) = "";
		(Bmult[22] => Cmult[4]) = "";
		(Bmult[23] => Cmult[4]) = "";
		(Bmult[24] => Cmult[4]) = "";
		(Bmult[25] => Cmult[4]) = "";
		(Bmult[26] => Cmult[4]) = "";
		(Bmult[27] => Cmult[4]) = "";
		(Bmult[28] => Cmult[4]) = "";
		(Bmult[29] => Cmult[4]) = "";
		(Bmult[30] => Cmult[4]) = "";
		(Bmult[31] => Cmult[4]) = "";		
		(Valid_mult[0] => Cmult[4]) = "";
		(Valid_mult[1] => Cmult[4]) = "";
		(sel_mul_32x32 => Cmult[4]) = "";
		(Amult[0]  => Cmult[5]) = "";
		(Amult[1]  => Cmult[5]) = "";
		(Amult[2]  => Cmult[5]) = "";
		(Amult[3]  => Cmult[5]) = "";
		(Amult[4]  => Cmult[5]) = "";
		(Amult[5]  => Cmult[5]) = "";
		(Amult[6]  => Cmult[5]) = "";
		(Amult[7]  => Cmult[5]) = "";
		(Amult[8]  => Cmult[5]) = "";
		(Amult[9]  => Cmult[5]) = "";
		(Amult[10] => Cmult[5]) = "";
		(Amult[11] => Cmult[5]) = "";
		(Amult[12] => Cmult[5]) = "";
		(Amult[13] => Cmult[5]) = "";
		(Amult[14] => Cmult[5]) = "";
		(Amult[15] => Cmult[5]) = "";
		(Amult[16] => Cmult[5]) = "";
		(Amult[17] => Cmult[5]) = "";
		(Amult[18] => Cmult[5]) = "";
		(Amult[19] => Cmult[5]) = "";
		(Amult[20] => Cmult[5]) = "";
		(Amult[21] => Cmult[5]) = "";
		(Amult[22] => Cmult[5]) = "";
		(Amult[23] => Cmult[5]) = "";
		(Amult[24] => Cmult[5]) = "";
		(Amult[25] => Cmult[5]) = "";
		(Amult[26] => Cmult[5]) = "";
		(Amult[27] => Cmult[5]) = "";
		(Amult[28] => Cmult[5]) = "";
		(Amult[29] => Cmult[5]) = "";
		(Amult[30] => Cmult[5]) = "";
		(Amult[31] => Cmult[5]) = "";
		(Bmult[0]  => Cmult[5]) = "";
		(Bmult[1]  => Cmult[5]) = "";
		(Bmult[2]  => Cmult[5]) = "";
		(Bmult[3]  => Cmult[5]) = "";
		(Bmult[4]  => Cmult[5]) = "";
		(Bmult[5]  => Cmult[5]) = "";
		(Bmult[6]  => Cmult[5]) = "";
		(Bmult[7]  => Cmult[5]) = "";
		(Bmult[8]  => Cmult[5]) = "";
		(Bmult[9]  => Cmult[5]) = "";
		(Bmult[10] => Cmult[5]) = "";
		(Bmult[11] => Cmult[5]) = "";
		(Bmult[12] => Cmult[5]) = "";
		(Bmult[13] => Cmult[5]) = "";
		(Bmult[14] => Cmult[5]) = "";
		(Bmult[15] => Cmult[5]) = "";
		(Bmult[16] => Cmult[5]) = "";
		(Bmult[17] => Cmult[5]) = "";
		(Bmult[18] => Cmult[5]) = "";
		(Bmult[19] => Cmult[5]) = "";
		(Bmult[20] => Cmult[5]) = "";
		(Bmult[21] => Cmult[5]) = "";
		(Bmult[22] => Cmult[5]) = "";
		(Bmult[23] => Cmult[5]) = "";
		(Bmult[24] => Cmult[5]) = "";
		(Bmult[25] => Cmult[5]) = "";
		(Bmult[26] => Cmult[5]) = "";
		(Bmult[27] => Cmult[5]) = "";
		(Bmult[28] => Cmult[5]) = "";
		(Bmult[29] => Cmult[5]) = "";
		(Bmult[30] => Cmult[5]) = "";
		(Bmult[31] => Cmult[5]) = "";		
		(Valid_mult[0] => Cmult[5]) = "";
		(Valid_mult[1] => Cmult[5]) = "";
		(sel_mul_32x32 => Cmult[5]) = "";
		(Amult[0]  => Cmult[6]) = "";
		(Amult[1]  => Cmult[6]) = "";
		(Amult[2]  => Cmult[6]) = "";
		(Amult[3]  => Cmult[6]) = "";
		(Amult[4]  => Cmult[6]) = "";
		(Amult[5]  => Cmult[6]) = "";
		(Amult[6]  => Cmult[6]) = "";
		(Amult[7]  => Cmult[6]) = "";
		(Amult[8]  => Cmult[6]) = "";
		(Amult[9]  => Cmult[6]) = "";
		(Amult[10] => Cmult[6]) = "";
		(Amult[11] => Cmult[6]) = "";
		(Amult[12] => Cmult[6]) = "";
		(Amult[13] => Cmult[6]) = "";
		(Amult[14] => Cmult[6]) = "";
		(Amult[15] => Cmult[6]) = "";
		(Amult[16] => Cmult[6]) = "";
		(Amult[17] => Cmult[6]) = "";
		(Amult[18] => Cmult[6]) = "";
		(Amult[19] => Cmult[6]) = "";
		(Amult[20] => Cmult[6]) = "";
		(Amult[21] => Cmult[6]) = "";
		(Amult[22] => Cmult[6]) = "";
		(Amult[23] => Cmult[6]) = "";
		(Amult[24] => Cmult[6]) = "";
		(Amult[25] => Cmult[6]) = "";
		(Amult[26] => Cmult[6]) = "";
		(Amult[27] => Cmult[6]) = "";
		(Amult[28] => Cmult[6]) = "";
		(Amult[29] => Cmult[6]) = "";
		(Amult[30] => Cmult[6]) = "";
		(Amult[31] => Cmult[6]) = "";
		(Bmult[0]  => Cmult[6]) = "";
		(Bmult[1]  => Cmult[6]) = "";
		(Bmult[2]  => Cmult[6]) = "";
		(Bmult[3]  => Cmult[6]) = "";
		(Bmult[4]  => Cmult[6]) = "";
		(Bmult[5]  => Cmult[6]) = "";
		(Bmult[6]  => Cmult[6]) = "";
		(Bmult[7]  => Cmult[6]) = "";
		(Bmult[8]  => Cmult[6]) = "";
		(Bmult[9]  => Cmult[6]) = "";
		(Bmult[10] => Cmult[6]) = "";
		(Bmult[11] => Cmult[6]) = "";
		(Bmult[12] => Cmult[6]) = "";
		(Bmult[13] => Cmult[6]) = "";
		(Bmult[14] => Cmult[6]) = "";
		(Bmult[15] => Cmult[6]) = "";
		(Bmult[16] => Cmult[6]) = "";
		(Bmult[17] => Cmult[6]) = "";
		(Bmult[18] => Cmult[6]) = "";
		(Bmult[19] => Cmult[6]) = "";
		(Bmult[20] => Cmult[6]) = "";
		(Bmult[21] => Cmult[6]) = "";
		(Bmult[22] => Cmult[6]) = "";
		(Bmult[23] => Cmult[6]) = "";
		(Bmult[24] => Cmult[6]) = "";
		(Bmult[25] => Cmult[6]) = "";
		(Bmult[26] => Cmult[6]) = "";
		(Bmult[27] => Cmult[6]) = "";
		(Bmult[28] => Cmult[6]) = "";
		(Bmult[29] => Cmult[6]) = "";
		(Bmult[30] => Cmult[6]) = "";
		(Bmult[31] => Cmult[6]) = "";		
		(Valid_mult[0] => Cmult[6]) = "";
		(Valid_mult[1] => Cmult[6]) = "";
		(sel_mul_32x32 => Cmult[6]) = "";
		(Amult[0]  => Cmult[7]) = "";
		(Amult[1]  => Cmult[7]) = "";
		(Amult[2]  => Cmult[7]) = "";
		(Amult[3]  => Cmult[7]) = "";
		(Amult[4]  => Cmult[7]) = "";
		(Amult[5]  => Cmult[7]) = "";
		(Amult[6]  => Cmult[7]) = "";
		(Amult[7]  => Cmult[7]) = "";
		(Amult[8]  => Cmult[7]) = "";
		(Amult[9]  => Cmult[7]) = "";
		(Amult[10] => Cmult[7]) = "";
		(Amult[11] => Cmult[7]) = "";
		(Amult[12] => Cmult[7]) = "";
		(Amult[13] => Cmult[7]) = "";
		(Amult[14] => Cmult[7]) = "";
		(Amult[15] => Cmult[7]) = "";
		(Amult[16] => Cmult[7]) = "";
		(Amult[17] => Cmult[7]) = "";
		(Amult[18] => Cmult[7]) = "";
		(Amult[19] => Cmult[7]) = "";
		(Amult[20] => Cmult[7]) = "";
		(Amult[21] => Cmult[7]) = "";
		(Amult[22] => Cmult[7]) = "";
		(Amult[23] => Cmult[7]) = "";
		(Amult[24] => Cmult[7]) = "";
		(Amult[25] => Cmult[7]) = "";
		(Amult[26] => Cmult[7]) = "";
		(Amult[27] => Cmult[7]) = "";
		(Amult[28] => Cmult[7]) = "";
		(Amult[29] => Cmult[7]) = "";
		(Amult[30] => Cmult[7]) = "";
		(Amult[31] => Cmult[7]) = "";
		(Bmult[0]  => Cmult[7]) = "";
		(Bmult[1]  => Cmult[7]) = "";
		(Bmult[2]  => Cmult[7]) = "";
		(Bmult[3]  => Cmult[7]) = "";
		(Bmult[4]  => Cmult[7]) = "";
		(Bmult[5]  => Cmult[7]) = "";
		(Bmult[6]  => Cmult[7]) = "";
		(Bmult[7]  => Cmult[7]) = "";
		(Bmult[8]  => Cmult[7]) = "";
		(Bmult[9]  => Cmult[7]) = "";
		(Bmult[10] => Cmult[7]) = "";
		(Bmult[11] => Cmult[7]) = "";
		(Bmult[12] => Cmult[7]) = "";
		(Bmult[13] => Cmult[7]) = "";
		(Bmult[14] => Cmult[7]) = "";
		(Bmult[15] => Cmult[7]) = "";
		(Bmult[16] => Cmult[7]) = "";
		(Bmult[17] => Cmult[7]) = "";
		(Bmult[18] => Cmult[7]) = "";
		(Bmult[19] => Cmult[7]) = "";
		(Bmult[20] => Cmult[7]) = "";
		(Bmult[21] => Cmult[7]) = "";
		(Bmult[22] => Cmult[7]) = "";
		(Bmult[23] => Cmult[7]) = "";
		(Bmult[24] => Cmult[7]) = "";
		(Bmult[25] => Cmult[7]) = "";
		(Bmult[26] => Cmult[7]) = "";
		(Bmult[27] => Cmult[7]) = "";
		(Bmult[28] => Cmult[7]) = "";
		(Bmult[29] => Cmult[7]) = "";
		(Bmult[30] => Cmult[7]) = "";
		(Bmult[31] => Cmult[7]) = "";		
		(Valid_mult[0] => Cmult[7]) = "";
		(Valid_mult[1] => Cmult[7]) = "";
		(sel_mul_32x32 => Cmult[7]) = "";
		(Amult[0]  => Cmult[8]) = "";
		(Amult[1]  => Cmult[8]) = "";
		(Amult[2]  => Cmult[8]) = "";
		(Amult[3]  => Cmult[8]) = "";
		(Amult[4]  => Cmult[8]) = "";
		(Amult[5]  => Cmult[8]) = "";
		(Amult[6]  => Cmult[8]) = "";
		(Amult[7]  => Cmult[8]) = "";
		(Amult[8]  => Cmult[8]) = "";
		(Amult[9]  => Cmult[8]) = "";
		(Amult[10] => Cmult[8]) = "";
		(Amult[11] => Cmult[8]) = "";
		(Amult[12] => Cmult[8]) = "";
		(Amult[13] => Cmult[8]) = "";
		(Amult[14] => Cmult[8]) = "";
		(Amult[15] => Cmult[8]) = "";
		(Amult[16] => Cmult[8]) = "";
		(Amult[17] => Cmult[8]) = "";
		(Amult[18] => Cmult[8]) = "";
		(Amult[19] => Cmult[8]) = "";
		(Amult[20] => Cmult[8]) = "";
		(Amult[21] => Cmult[8]) = "";
		(Amult[22] => Cmult[8]) = "";
		(Amult[23] => Cmult[8]) = "";
		(Amult[24] => Cmult[8]) = "";
		(Amult[25] => Cmult[8]) = "";
		(Amult[26] => Cmult[8]) = "";
		(Amult[27] => Cmult[8]) = "";
		(Amult[28] => Cmult[8]) = "";
		(Amult[29] => Cmult[8]) = "";
		(Amult[30] => Cmult[8]) = "";
		(Amult[31] => Cmult[8]) = "";
		(Bmult[0]  => Cmult[8]) = "";
		(Bmult[1]  => Cmult[8]) = "";
		(Bmult[2]  => Cmult[8]) = "";
		(Bmult[3]  => Cmult[8]) = "";
		(Bmult[4]  => Cmult[8]) = "";
		(Bmult[5]  => Cmult[8]) = "";
		(Bmult[6]  => Cmult[8]) = "";
		(Bmult[7]  => Cmult[8]) = "";
		(Bmult[8]  => Cmult[8]) = "";
		(Bmult[9]  => Cmult[8]) = "";
		(Bmult[10] => Cmult[8]) = "";
		(Bmult[11] => Cmult[8]) = "";
		(Bmult[12] => Cmult[8]) = "";
		(Bmult[13] => Cmult[8]) = "";
		(Bmult[14] => Cmult[8]) = "";
		(Bmult[15] => Cmult[8]) = "";
		(Bmult[16] => Cmult[8]) = "";
		(Bmult[17] => Cmult[8]) = "";
		(Bmult[18] => Cmult[8]) = "";
		(Bmult[19] => Cmult[8]) = "";
		(Bmult[20] => Cmult[8]) = "";
		(Bmult[21] => Cmult[8]) = "";
		(Bmult[22] => Cmult[8]) = "";
		(Bmult[23] => Cmult[8]) = "";
		(Bmult[24] => Cmult[8]) = "";
		(Bmult[25] => Cmult[8]) = "";
		(Bmult[26] => Cmult[8]) = "";
		(Bmult[27] => Cmult[8]) = "";
		(Bmult[28] => Cmult[8]) = "";
		(Bmult[29] => Cmult[8]) = "";
		(Bmult[30] => Cmult[8]) = "";
		(Bmult[31] => Cmult[8]) = "";		
		(Valid_mult[0] => Cmult[8]) = "";
		(Valid_mult[1] => Cmult[8]) = "";
		(sel_mul_32x32 => Cmult[8]) = "";	
		(Amult[0]  => Cmult[9]) = "";
		(Amult[1]  => Cmult[9]) = "";
		(Amult[2]  => Cmult[9]) = "";
		(Amult[3]  => Cmult[9]) = "";
		(Amult[4]  => Cmult[9]) = "";
		(Amult[5]  => Cmult[9]) = "";
		(Amult[6]  => Cmult[9]) = "";
		(Amult[7]  => Cmult[9]) = "";
		(Amult[8]  => Cmult[9]) = "";
		(Amult[9]  => Cmult[9]) = "";
		(Amult[10] => Cmult[9]) = "";
		(Amult[11] => Cmult[9]) = "";
		(Amult[12] => Cmult[9]) = "";
		(Amult[13] => Cmult[9]) = "";
		(Amult[14] => Cmult[9]) = "";
		(Amult[15] => Cmult[9]) = "";
		(Amult[16] => Cmult[9]) = "";
		(Amult[17] => Cmult[9]) = "";
		(Amult[18] => Cmult[9]) = "";
		(Amult[19] => Cmult[9]) = "";
		(Amult[20] => Cmult[9]) = "";
		(Amult[21] => Cmult[9]) = "";
		(Amult[22] => Cmult[9]) = "";
		(Amult[23] => Cmult[9]) = "";
		(Amult[24] => Cmult[9]) = "";
		(Amult[25] => Cmult[9]) = "";
		(Amult[26] => Cmult[9]) = "";
		(Amult[27] => Cmult[9]) = "";
		(Amult[28] => Cmult[9]) = "";
		(Amult[29] => Cmult[9]) = "";
		(Amult[30] => Cmult[9]) = "";
		(Amult[31] => Cmult[9]) = "";
		(Bmult[0]  => Cmult[9]) = "";
		(Bmult[1]  => Cmult[9]) = "";
		(Bmult[2]  => Cmult[9]) = "";
		(Bmult[3]  => Cmult[9]) = "";
		(Bmult[4]  => Cmult[9]) = "";
		(Bmult[5]  => Cmult[9]) = "";
		(Bmult[6]  => Cmult[9]) = "";
		(Bmult[7]  => Cmult[9]) = "";
		(Bmult[8]  => Cmult[9]) = "";
		(Bmult[9]  => Cmult[9]) = "";
		(Bmult[10] => Cmult[9]) = "";
		(Bmult[11] => Cmult[9]) = "";
		(Bmult[12] => Cmult[9]) = "";
		(Bmult[13] => Cmult[9]) = "";
		(Bmult[14] => Cmult[9]) = "";
		(Bmult[15] => Cmult[9]) = "";
		(Bmult[16] => Cmult[9]) = "";
		(Bmult[17] => Cmult[9]) = "";
		(Bmult[18] => Cmult[9]) = "";
		(Bmult[19] => Cmult[9]) = "";
		(Bmult[20] => Cmult[9]) = "";
		(Bmult[21] => Cmult[9]) = "";
		(Bmult[22] => Cmult[9]) = "";
		(Bmult[23] => Cmult[9]) = "";
		(Bmult[24] => Cmult[9]) = "";
		(Bmult[25] => Cmult[9]) = "";
		(Bmult[26] => Cmult[9]) = "";
		(Bmult[27] => Cmult[9]) = "";
		(Bmult[28] => Cmult[9]) = "";
		(Bmult[29] => Cmult[9]) = "";
		(Bmult[30] => Cmult[9]) = "";
		(Bmult[31] => Cmult[9]) = "";		
		(Valid_mult[0] => Cmult[9]) = "";
		(Valid_mult[1] => Cmult[9]) = "";
		(sel_mul_32x32 => Cmult[9]) = "";	
		(Amult[0]  => Cmult[10]) = "";
		(Amult[1]  => Cmult[10]) = "";
		(Amult[2]  => Cmult[10]) = "";
		(Amult[3]  => Cmult[10]) = "";
		(Amult[4]  => Cmult[10]) = "";
		(Amult[5]  => Cmult[10]) = "";
		(Amult[6]  => Cmult[10]) = "";
		(Amult[7]  => Cmult[10]) = "";
		(Amult[8]  => Cmult[10]) = "";
		(Amult[9]  => Cmult[10]) = "";
		(Amult[10] => Cmult[10]) = "";
		(Amult[11] => Cmult[10]) = "";
		(Amult[12] => Cmult[10]) = "";
		(Amult[13] => Cmult[10]) = "";
		(Amult[14] => Cmult[10]) = "";
		(Amult[15] => Cmult[10]) = "";
		(Amult[16] => Cmult[10]) = "";
		(Amult[17] => Cmult[10]) = "";
		(Amult[18] => Cmult[10]) = "";
		(Amult[19] => Cmult[10]) = "";
		(Amult[20] => Cmult[10]) = "";
		(Amult[21] => Cmult[10]) = "";
		(Amult[22] => Cmult[10]) = "";
		(Amult[23] => Cmult[10]) = "";
		(Amult[24] => Cmult[10]) = "";
		(Amult[25] => Cmult[10]) = "";
		(Amult[26] => Cmult[10]) = "";
		(Amult[27] => Cmult[10]) = "";
		(Amult[28] => Cmult[10]) = "";
		(Amult[29] => Cmult[10]) = "";
		(Amult[30] => Cmult[10]) = "";
		(Amult[31] => Cmult[10]) = "";
		(Bmult[0]  => Cmult[10]) = "";
		(Bmult[1]  => Cmult[10]) = "";
		(Bmult[2]  => Cmult[10]) = "";
		(Bmult[3]  => Cmult[10]) = "";
		(Bmult[4]  => Cmult[10]) = "";
		(Bmult[5]  => Cmult[10]) = "";
		(Bmult[6]  => Cmult[10]) = "";
		(Bmult[7]  => Cmult[10]) = "";
		(Bmult[8]  => Cmult[10]) = "";
		(Bmult[9]  => Cmult[10]) = "";
		(Bmult[10] => Cmult[10]) = "";
		(Bmult[11] => Cmult[10]) = "";
		(Bmult[12] => Cmult[10]) = "";
		(Bmult[13] => Cmult[10]) = "";
		(Bmult[14] => Cmult[10]) = "";
		(Bmult[15] => Cmult[10]) = "";
		(Bmult[16] => Cmult[10]) = "";
		(Bmult[17] => Cmult[10]) = "";
		(Bmult[18] => Cmult[10]) = "";
		(Bmult[19] => Cmult[10]) = "";
		(Bmult[20] => Cmult[10]) = "";
		(Bmult[21] => Cmult[10]) = "";
		(Bmult[22] => Cmult[10]) = "";
		(Bmult[23] => Cmult[10]) = "";
		(Bmult[24] => Cmult[10]) = "";
		(Bmult[25] => Cmult[10]) = "";
		(Bmult[26] => Cmult[10]) = "";
		(Bmult[27] => Cmult[10]) = "";
		(Bmult[28] => Cmult[10]) = "";
		(Bmult[29] => Cmult[10]) = "";
		(Bmult[30] => Cmult[10]) = "";
		(Bmult[31] => Cmult[10]) = "";		
		(Valid_mult[0] => Cmult[10]) = "";
		(Valid_mult[1] => Cmult[10]) = "";
		(sel_mul_32x32 => Cmult[10]) = "";
		(Amult[0]  => Cmult[11]) = "";
		(Amult[1]  => Cmult[11]) = "";
		(Amult[2]  => Cmult[11]) = "";
		(Amult[3]  => Cmult[11]) = "";
		(Amult[4]  => Cmult[11]) = "";
		(Amult[5]  => Cmult[11]) = "";
		(Amult[6]  => Cmult[11]) = "";
		(Amult[7]  => Cmult[11]) = "";
		(Amult[8]  => Cmult[11]) = "";
		(Amult[9]  => Cmult[11]) = "";
		(Amult[10] => Cmult[11]) = "";
		(Amult[11] => Cmult[11]) = "";
		(Amult[12] => Cmult[11]) = "";
		(Amult[13] => Cmult[11]) = "";
		(Amult[14] => Cmult[11]) = "";
		(Amult[15] => Cmult[11]) = "";
		(Amult[16] => Cmult[11]) = "";
		(Amult[17] => Cmult[11]) = "";
		(Amult[18] => Cmult[11]) = "";
		(Amult[19] => Cmult[11]) = "";
		(Amult[20] => Cmult[11]) = "";
		(Amult[21] => Cmult[11]) = "";
		(Amult[22] => Cmult[11]) = "";
		(Amult[23] => Cmult[11]) = "";
		(Amult[24] => Cmult[11]) = "";
		(Amult[25] => Cmult[11]) = "";
		(Amult[26] => Cmult[11]) = "";
		(Amult[27] => Cmult[11]) = "";
		(Amult[28] => Cmult[11]) = "";
		(Amult[29] => Cmult[11]) = "";
		(Amult[30] => Cmult[11]) = "";
		(Amult[31] => Cmult[11]) = "";
		(Bmult[0]  => Cmult[11]) = "";
		(Bmult[1]  => Cmult[11]) = "";
		(Bmult[2]  => Cmult[11]) = "";
		(Bmult[3]  => Cmult[11]) = "";
		(Bmult[4]  => Cmult[11]) = "";
		(Bmult[5]  => Cmult[11]) = "";
		(Bmult[6]  => Cmult[11]) = "";
		(Bmult[7]  => Cmult[11]) = "";
		(Bmult[8]  => Cmult[11]) = "";
		(Bmult[9]  => Cmult[11]) = "";
		(Bmult[10] => Cmult[11]) = "";
		(Bmult[11] => Cmult[11]) = "";
		(Bmult[12] => Cmult[11]) = "";
		(Bmult[13] => Cmult[11]) = "";
		(Bmult[14] => Cmult[11]) = "";
		(Bmult[15] => Cmult[11]) = "";
		(Bmult[16] => Cmult[11]) = "";
		(Bmult[17] => Cmult[11]) = "";
		(Bmult[18] => Cmult[11]) = "";
		(Bmult[19] => Cmult[11]) = "";
		(Bmult[20] => Cmult[11]) = "";
		(Bmult[21] => Cmult[11]) = "";
		(Bmult[22] => Cmult[11]) = "";
		(Bmult[23] => Cmult[11]) = "";
		(Bmult[24] => Cmult[11]) = "";
		(Bmult[25] => Cmult[11]) = "";
		(Bmult[26] => Cmult[11]) = "";
		(Bmult[27] => Cmult[11]) = "";
		(Bmult[28] => Cmult[11]) = "";
		(Bmult[29] => Cmult[11]) = "";
		(Bmult[30] => Cmult[11]) = "";
		(Bmult[31] => Cmult[11]) = "";		
		(Valid_mult[0] => Cmult[11]) = "";
		(Valid_mult[1] => Cmult[11]) = "";
		(sel_mul_32x32 => Cmult[11]) = "";
		(Amult[0]  => Cmult[12]) = "";
		(Amult[1]  => Cmult[12]) = "";
		(Amult[2]  => Cmult[12]) = "";
		(Amult[3]  => Cmult[12]) = "";
		(Amult[4]  => Cmult[12]) = "";
		(Amult[5]  => Cmult[12]) = "";
		(Amult[6]  => Cmult[12]) = "";
		(Amult[7]  => Cmult[12]) = "";
		(Amult[8]  => Cmult[12]) = "";
		(Amult[9]  => Cmult[12]) = "";
		(Amult[10] => Cmult[12]) = "";
		(Amult[11] => Cmult[12]) = "";
		(Amult[12] => Cmult[12]) = "";
		(Amult[13] => Cmult[12]) = "";
		(Amult[14] => Cmult[12]) = "";
		(Amult[15] => Cmult[12]) = "";
		(Amult[16] => Cmult[12]) = "";
		(Amult[17] => Cmult[12]) = "";
		(Amult[18] => Cmult[12]) = "";
		(Amult[19] => Cmult[12]) = "";
		(Amult[20] => Cmult[12]) = "";
		(Amult[21] => Cmult[12]) = "";
		(Amult[22] => Cmult[12]) = "";
		(Amult[23] => Cmult[12]) = "";
		(Amult[24] => Cmult[12]) = "";
		(Amult[25] => Cmult[12]) = "";
		(Amult[26] => Cmult[12]) = "";
		(Amult[27] => Cmult[12]) = "";
		(Amult[28] => Cmult[12]) = "";
		(Amult[29] => Cmult[12]) = "";
		(Amult[30] => Cmult[12]) = "";
		(Amult[31] => Cmult[12]) = "";
		(Bmult[0]  => Cmult[12]) = "";
		(Bmult[1]  => Cmult[12]) = "";
		(Bmult[2]  => Cmult[12]) = "";
		(Bmult[3]  => Cmult[12]) = "";
		(Bmult[4]  => Cmult[12]) = "";
		(Bmult[5]  => Cmult[12]) = "";
		(Bmult[6]  => Cmult[12]) = "";
		(Bmult[7]  => Cmult[12]) = "";
		(Bmult[8]  => Cmult[12]) = "";
		(Bmult[9]  => Cmult[12]) = "";
		(Bmult[10] => Cmult[12]) = "";
		(Bmult[11] => Cmult[12]) = "";
		(Bmult[12] => Cmult[12]) = "";
		(Bmult[13] => Cmult[12]) = "";
		(Bmult[14] => Cmult[12]) = "";
		(Bmult[15] => Cmult[12]) = "";
		(Bmult[16] => Cmult[12]) = "";
		(Bmult[17] => Cmult[12]) = "";
		(Bmult[18] => Cmult[12]) = "";
		(Bmult[19] => Cmult[12]) = "";
		(Bmult[20] => Cmult[12]) = "";
		(Bmult[21] => Cmult[12]) = "";
		(Bmult[22] => Cmult[12]) = "";
		(Bmult[23] => Cmult[12]) = "";
		(Bmult[24] => Cmult[12]) = "";
		(Bmult[25] => Cmult[12]) = "";
		(Bmult[26] => Cmult[12]) = "";
		(Bmult[27] => Cmult[12]) = "";
		(Bmult[28] => Cmult[12]) = "";
		(Bmult[29] => Cmult[12]) = "";
		(Bmult[30] => Cmult[12]) = "";
		(Bmult[31] => Cmult[12]) = "";		
		(Valid_mult[0] => Cmult[12]) = "";
		(Valid_mult[1] => Cmult[12]) = "";
		(sel_mul_32x32 => Cmult[12]) = "";
		(Amult[0]  => Cmult[13]) = "";
		(Amult[1]  => Cmult[13]) = "";
		(Amult[2]  => Cmult[13]) = "";
		(Amult[3]  => Cmult[13]) = "";
		(Amult[4]  => Cmult[13]) = "";
		(Amult[5]  => Cmult[13]) = "";
		(Amult[6]  => Cmult[13]) = "";
		(Amult[7]  => Cmult[13]) = "";
		(Amult[8]  => Cmult[13]) = "";
		(Amult[9]  => Cmult[13]) = "";
		(Amult[10] => Cmult[13]) = "";
		(Amult[11] => Cmult[13]) = "";
		(Amult[12] => Cmult[13]) = "";
		(Amult[13] => Cmult[13]) = "";
		(Amult[14] => Cmult[13]) = "";
		(Amult[15] => Cmult[13]) = "";
		(Amult[16] => Cmult[13]) = "";
		(Amult[17] => Cmult[13]) = "";
		(Amult[18] => Cmult[13]) = "";
		(Amult[19] => Cmult[13]) = "";
		(Amult[20] => Cmult[13]) = "";
		(Amult[21] => Cmult[13]) = "";
		(Amult[22] => Cmult[13]) = "";
		(Amult[23] => Cmult[13]) = "";
		(Amult[24] => Cmult[13]) = "";
		(Amult[25] => Cmult[13]) = "";
		(Amult[26] => Cmult[13]) = "";
		(Amult[27] => Cmult[13]) = "";
		(Amult[28] => Cmult[13]) = "";
		(Amult[29] => Cmult[13]) = "";
		(Amult[30] => Cmult[13]) = "";
		(Amult[31] => Cmult[13]) = "";
		(Bmult[0]  => Cmult[13]) = "";
		(Bmult[1]  => Cmult[13]) = "";
		(Bmult[2]  => Cmult[13]) = "";
		(Bmult[3]  => Cmult[13]) = "";
		(Bmult[4]  => Cmult[13]) = "";
		(Bmult[5]  => Cmult[13]) = "";
		(Bmult[6]  => Cmult[13]) = "";
		(Bmult[7]  => Cmult[13]) = "";
		(Bmult[8]  => Cmult[13]) = "";
		(Bmult[9]  => Cmult[13]) = "";
		(Bmult[10] => Cmult[13]) = "";
		(Bmult[11] => Cmult[13]) = "";
		(Bmult[12] => Cmult[13]) = "";
		(Bmult[13] => Cmult[13]) = "";
		(Bmult[14] => Cmult[13]) = "";
		(Bmult[15] => Cmult[13]) = "";
		(Bmult[16] => Cmult[13]) = "";
		(Bmult[17] => Cmult[13]) = "";
		(Bmult[18] => Cmult[13]) = "";
		(Bmult[19] => Cmult[13]) = "";
		(Bmult[20] => Cmult[13]) = "";
		(Bmult[21] => Cmult[13]) = "";
		(Bmult[22] => Cmult[13]) = "";
		(Bmult[23] => Cmult[13]) = "";
		(Bmult[24] => Cmult[13]) = "";
		(Bmult[25] => Cmult[13]) = "";
		(Bmult[26] => Cmult[13]) = "";
		(Bmult[27] => Cmult[13]) = "";
		(Bmult[28] => Cmult[13]) = "";
		(Bmult[29] => Cmult[13]) = "";
		(Bmult[30] => Cmult[13]) = "";
		(Bmult[31] => Cmult[13]) = "";		
		(Valid_mult[0] => Cmult[13]) = "";
		(Valid_mult[1] => Cmult[13]) = "";
		(sel_mul_32x32 => Cmult[13]) = "";
		(Amult[0]  => Cmult[14]) = "";
		(Amult[1]  => Cmult[14]) = "";
		(Amult[2]  => Cmult[14]) = "";
		(Amult[3]  => Cmult[14]) = "";
		(Amult[4]  => Cmult[14]) = "";
		(Amult[5]  => Cmult[14]) = "";
		(Amult[6]  => Cmult[14]) = "";
		(Amult[7]  => Cmult[14]) = "";
		(Amult[8]  => Cmult[14]) = "";
		(Amult[9]  => Cmult[14]) = "";
		(Amult[10] => Cmult[14]) = "";
		(Amult[11] => Cmult[14]) = "";
		(Amult[12] => Cmult[14]) = "";
		(Amult[13] => Cmult[14]) = "";
		(Amult[14] => Cmult[14]) = "";
		(Amult[15] => Cmult[14]) = "";
		(Amult[16] => Cmult[14]) = "";
		(Amult[17] => Cmult[14]) = "";
		(Amult[18] => Cmult[14]) = "";
		(Amult[19] => Cmult[14]) = "";
		(Amult[20] => Cmult[14]) = "";
		(Amult[21] => Cmult[14]) = "";
		(Amult[22] => Cmult[14]) = "";
		(Amult[23] => Cmult[14]) = "";
		(Amult[24] => Cmult[14]) = "";
		(Amult[25] => Cmult[14]) = "";
		(Amult[26] => Cmult[14]) = "";
		(Amult[27] => Cmult[14]) = "";
		(Amult[28] => Cmult[14]) = "";
		(Amult[29] => Cmult[14]) = "";
		(Amult[30] => Cmult[14]) = "";
		(Amult[31] => Cmult[14]) = "";
		(Bmult[0]  => Cmult[14]) = "";
		(Bmult[1]  => Cmult[14]) = "";
		(Bmult[2]  => Cmult[14]) = "";
		(Bmult[3]  => Cmult[14]) = "";
		(Bmult[4]  => Cmult[14]) = "";
		(Bmult[5]  => Cmult[14]) = "";
		(Bmult[6]  => Cmult[14]) = "";
		(Bmult[7]  => Cmult[14]) = "";
		(Bmult[8]  => Cmult[14]) = "";
		(Bmult[9]  => Cmult[14]) = "";
		(Bmult[10] => Cmult[14]) = "";
		(Bmult[11] => Cmult[14]) = "";
		(Bmult[12] => Cmult[14]) = "";
		(Bmult[13] => Cmult[14]) = "";
		(Bmult[14] => Cmult[14]) = "";
		(Bmult[15] => Cmult[14]) = "";
		(Bmult[16] => Cmult[14]) = "";
		(Bmult[17] => Cmult[14]) = "";
		(Bmult[18] => Cmult[14]) = "";
		(Bmult[19] => Cmult[14]) = "";
		(Bmult[20] => Cmult[14]) = "";
		(Bmult[21] => Cmult[14]) = "";
		(Bmult[22] => Cmult[14]) = "";
		(Bmult[23] => Cmult[14]) = "";
		(Bmult[24] => Cmult[14]) = "";
		(Bmult[25] => Cmult[14]) = "";
		(Bmult[26] => Cmult[14]) = "";
		(Bmult[27] => Cmult[14]) = "";
		(Bmult[28] => Cmult[14]) = "";
		(Bmult[29] => Cmult[14]) = "";
		(Bmult[30] => Cmult[14]) = "";
		(Bmult[31] => Cmult[14]) = "";		
		(Valid_mult[0] => Cmult[14]) = "";
		(Valid_mult[1] => Cmult[14]) = "";
		(sel_mul_32x32 => Cmult[14]) = "";
		(Amult[0]  => Cmult[15]) = "";
		(Amult[1]  => Cmult[15]) = "";
		(Amult[2]  => Cmult[15]) = "";
		(Amult[3]  => Cmult[15]) = "";
		(Amult[4]  => Cmult[15]) = "";
		(Amult[5]  => Cmult[15]) = "";
		(Amult[6]  => Cmult[15]) = "";
		(Amult[7]  => Cmult[15]) = "";
		(Amult[8]  => Cmult[15]) = "";
		(Amult[9]  => Cmult[15]) = "";
		(Amult[10] => Cmult[15]) = "";
		(Amult[11] => Cmult[15]) = "";
		(Amult[12] => Cmult[15]) = "";
		(Amult[13] => Cmult[15]) = "";
		(Amult[14] => Cmult[15]) = "";
		(Amult[15] => Cmult[15]) = "";
		(Amult[16] => Cmult[15]) = "";
		(Amult[17] => Cmult[15]) = "";
		(Amult[18] => Cmult[15]) = "";
		(Amult[19] => Cmult[15]) = "";
		(Amult[20] => Cmult[15]) = "";
		(Amult[21] => Cmult[15]) = "";
		(Amult[22] => Cmult[15]) = "";
		(Amult[23] => Cmult[15]) = "";
		(Amult[24] => Cmult[15]) = "";
		(Amult[25] => Cmult[15]) = "";
		(Amult[26] => Cmult[15]) = "";
		(Amult[27] => Cmult[15]) = "";
		(Amult[28] => Cmult[15]) = "";
		(Amult[29] => Cmult[15]) = "";
		(Amult[30] => Cmult[15]) = "";
		(Amult[31] => Cmult[15]) = "";
		(Bmult[0]  => Cmult[15]) = "";
		(Bmult[1]  => Cmult[15]) = "";
		(Bmult[2]  => Cmult[15]) = "";
		(Bmult[3]  => Cmult[15]) = "";
		(Bmult[4]  => Cmult[15]) = "";
		(Bmult[5]  => Cmult[15]) = "";
		(Bmult[6]  => Cmult[15]) = "";
		(Bmult[7]  => Cmult[15]) = "";
		(Bmult[8]  => Cmult[15]) = "";
		(Bmult[9]  => Cmult[15]) = "";
		(Bmult[10] => Cmult[15]) = "";
		(Bmult[11] => Cmult[15]) = "";
		(Bmult[12] => Cmult[15]) = "";
		(Bmult[13] => Cmult[15]) = "";
		(Bmult[14] => Cmult[15]) = "";
		(Bmult[15] => Cmult[15]) = "";
		(Bmult[16] => Cmult[15]) = "";
		(Bmult[17] => Cmult[15]) = "";
		(Bmult[18] => Cmult[15]) = "";
		(Bmult[19] => Cmult[15]) = "";
		(Bmult[20] => Cmult[15]) = "";
		(Bmult[21] => Cmult[15]) = "";
		(Bmult[22] => Cmult[15]) = "";
		(Bmult[23] => Cmult[15]) = "";
		(Bmult[24] => Cmult[15]) = "";
		(Bmult[25] => Cmult[15]) = "";
		(Bmult[26] => Cmult[15]) = "";
		(Bmult[27] => Cmult[15]) = "";
		(Bmult[28] => Cmult[15]) = "";
		(Bmult[29] => Cmult[15]) = "";
		(Bmult[30] => Cmult[15]) = "";
		(Bmult[31] => Cmult[15]) = "";		
		(Valid_mult[0] => Cmult[15]) = "";
		(Valid_mult[1] => Cmult[15]) = "";
		(sel_mul_32x32 => Cmult[15]) = "";
		(Amult[0]  => Cmult[16]) = "";
		(Amult[1]  => Cmult[16]) = "";
		(Amult[2]  => Cmult[16]) = "";
		(Amult[3]  => Cmult[16]) = "";
		(Amult[4]  => Cmult[16]) = "";
		(Amult[5]  => Cmult[16]) = "";
		(Amult[6]  => Cmult[16]) = "";
		(Amult[7]  => Cmult[16]) = "";
		(Amult[8]  => Cmult[16]) = "";
		(Amult[9]  => Cmult[16]) = "";
		(Amult[10] => Cmult[16]) = "";
		(Amult[11] => Cmult[16]) = "";
		(Amult[12] => Cmult[16]) = "";
		(Amult[13] => Cmult[16]) = "";
		(Amult[14] => Cmult[16]) = "";
		(Amult[15] => Cmult[16]) = "";
		(Amult[16] => Cmult[16]) = "";
		(Amult[17] => Cmult[16]) = "";
		(Amult[18] => Cmult[16]) = "";
		(Amult[19] => Cmult[16]) = "";
		(Amult[20] => Cmult[16]) = "";
		(Amult[21] => Cmult[16]) = "";
		(Amult[22] => Cmult[16]) = "";
		(Amult[23] => Cmult[16]) = "";
		(Amult[24] => Cmult[16]) = "";
		(Amult[25] => Cmult[16]) = "";
		(Amult[26] => Cmult[16]) = "";
		(Amult[27] => Cmult[16]) = "";
		(Amult[28] => Cmult[16]) = "";
		(Amult[29] => Cmult[16]) = "";
		(Amult[30] => Cmult[16]) = "";
		(Amult[31] => Cmult[16]) = "";
		(Bmult[0]  => Cmult[16]) = "";
		(Bmult[1]  => Cmult[16]) = "";
		(Bmult[2]  => Cmult[16]) = "";
		(Bmult[3]  => Cmult[16]) = "";
		(Bmult[4]  => Cmult[16]) = "";
		(Bmult[5]  => Cmult[16]) = "";
		(Bmult[6]  => Cmult[16]) = "";
		(Bmult[7]  => Cmult[16]) = "";
		(Bmult[8]  => Cmult[16]) = "";
		(Bmult[9]  => Cmult[16]) = "";
		(Bmult[10] => Cmult[16]) = "";
		(Bmult[11] => Cmult[16]) = "";
		(Bmult[12] => Cmult[16]) = "";
		(Bmult[13] => Cmult[16]) = "";
		(Bmult[14] => Cmult[16]) = "";
		(Bmult[15] => Cmult[16]) = "";
		(Bmult[16] => Cmult[16]) = "";
		(Bmult[17] => Cmult[16]) = "";
		(Bmult[18] => Cmult[16]) = "";
		(Bmult[19] => Cmult[16]) = "";
		(Bmult[20] => Cmult[16]) = "";
		(Bmult[21] => Cmult[16]) = "";
		(Bmult[22] => Cmult[16]) = "";
		(Bmult[23] => Cmult[16]) = "";
		(Bmult[24] => Cmult[16]) = "";
		(Bmult[25] => Cmult[16]) = "";
		(Bmult[26] => Cmult[16]) = "";
		(Bmult[27] => Cmult[16]) = "";
		(Bmult[28] => Cmult[16]) = "";
		(Bmult[29] => Cmult[16]) = "";
		(Bmult[30] => Cmult[16]) = "";
		(Bmult[31] => Cmult[16]) = "";		
		(Valid_mult[0] => Cmult[16]) = "";
		(Valid_mult[1] => Cmult[16]) = "";
		(sel_mul_32x32 => Cmult[16]) = "";
		(Amult[0]  => Cmult[17]) = "";
		(Amult[1]  => Cmult[17]) = "";
		(Amult[2]  => Cmult[17]) = "";
		(Amult[3]  => Cmult[17]) = "";
		(Amult[4]  => Cmult[17]) = "";
		(Amult[5]  => Cmult[17]) = "";
		(Amult[6]  => Cmult[17]) = "";
		(Amult[7]  => Cmult[17]) = "";
		(Amult[8]  => Cmult[17]) = "";
		(Amult[9]  => Cmult[17]) = "";
		(Amult[10] => Cmult[17]) = "";
		(Amult[11] => Cmult[17]) = "";
		(Amult[12] => Cmult[17]) = "";
		(Amult[13] => Cmult[17]) = "";
		(Amult[14] => Cmult[17]) = "";
		(Amult[15] => Cmult[17]) = "";
		(Amult[16] => Cmult[17]) = "";
		(Amult[17] => Cmult[17]) = "";
		(Amult[18] => Cmult[17]) = "";
		(Amult[19] => Cmult[17]) = "";
		(Amult[20] => Cmult[17]) = "";
		(Amult[21] => Cmult[17]) = "";
		(Amult[22] => Cmult[17]) = "";
		(Amult[23] => Cmult[17]) = "";
		(Amult[24] => Cmult[17]) = "";
		(Amult[25] => Cmult[17]) = "";
		(Amult[26] => Cmult[17]) = "";
		(Amult[27] => Cmult[17]) = "";
		(Amult[28] => Cmult[17]) = "";
		(Amult[29] => Cmult[17]) = "";
		(Amult[30] => Cmult[17]) = "";
		(Amult[31] => Cmult[17]) = "";
		(Bmult[0]  => Cmult[17]) = "";
		(Bmult[1]  => Cmult[17]) = "";
		(Bmult[2]  => Cmult[17]) = "";
		(Bmult[3]  => Cmult[17]) = "";
		(Bmult[4]  => Cmult[17]) = "";
		(Bmult[5]  => Cmult[17]) = "";
		(Bmult[6]  => Cmult[17]) = "";
		(Bmult[7]  => Cmult[17]) = "";
		(Bmult[8]  => Cmult[17]) = "";
		(Bmult[9]  => Cmult[17]) = "";
		(Bmult[10] => Cmult[17]) = "";
		(Bmult[11] => Cmult[17]) = "";
		(Bmult[12] => Cmult[17]) = "";
		(Bmult[13] => Cmult[17]) = "";
		(Bmult[14] => Cmult[17]) = "";
		(Bmult[15] => Cmult[17]) = "";
		(Bmult[16] => Cmult[17]) = "";
		(Bmult[17] => Cmult[17]) = "";
		(Bmult[18] => Cmult[17]) = "";
		(Bmult[19] => Cmult[17]) = "";
		(Bmult[20] => Cmult[17]) = "";
		(Bmult[21] => Cmult[17]) = "";
		(Bmult[22] => Cmult[17]) = "";
		(Bmult[23] => Cmult[17]) = "";
		(Bmult[24] => Cmult[17]) = "";
		(Bmult[25] => Cmult[17]) = "";
		(Bmult[26] => Cmult[17]) = "";
		(Bmult[27] => Cmult[17]) = "";
		(Bmult[28] => Cmult[17]) = "";
		(Bmult[29] => Cmult[17]) = "";
		(Bmult[30] => Cmult[17]) = "";
		(Bmult[31] => Cmult[17]) = "";		
		(Valid_mult[0] => Cmult[17]) = "";
		(Valid_mult[1] => Cmult[17]) = "";
		(sel_mul_32x32 => Cmult[17]) = "";
		(Amult[0]  => Cmult[18]) = "";
		(Amult[1]  => Cmult[18]) = "";
		(Amult[2]  => Cmult[18]) = "";
		(Amult[3]  => Cmult[18]) = "";
		(Amult[4]  => Cmult[18]) = "";
		(Amult[5]  => Cmult[18]) = "";
		(Amult[6]  => Cmult[18]) = "";
		(Amult[7]  => Cmult[18]) = "";
		(Amult[8]  => Cmult[18]) = "";
		(Amult[9]  => Cmult[18]) = "";
		(Amult[10] => Cmult[18]) = "";
		(Amult[11] => Cmult[18]) = "";
		(Amult[12] => Cmult[18]) = "";
		(Amult[13] => Cmult[18]) = "";
		(Amult[14] => Cmult[18]) = "";
		(Amult[15] => Cmult[18]) = "";
		(Amult[16] => Cmult[18]) = "";
		(Amult[17] => Cmult[18]) = "";
		(Amult[18] => Cmult[18]) = "";
		(Amult[19] => Cmult[18]) = "";
		(Amult[20] => Cmult[18]) = "";
		(Amult[21] => Cmult[18]) = "";
		(Amult[22] => Cmult[18]) = "";
		(Amult[23] => Cmult[18]) = "";
		(Amult[24] => Cmult[18]) = "";
		(Amult[25] => Cmult[18]) = "";
		(Amult[26] => Cmult[18]) = "";
		(Amult[27] => Cmult[18]) = "";
		(Amult[28] => Cmult[18]) = "";
		(Amult[29] => Cmult[18]) = "";
		(Amult[30] => Cmult[18]) = "";
		(Amult[31] => Cmult[18]) = "";
		(Bmult[0]  => Cmult[18]) = "";
		(Bmult[1]  => Cmult[18]) = "";
		(Bmult[2]  => Cmult[18]) = "";
		(Bmult[3]  => Cmult[18]) = "";
		(Bmult[4]  => Cmult[18]) = "";
		(Bmult[5]  => Cmult[18]) = "";
		(Bmult[6]  => Cmult[18]) = "";
		(Bmult[7]  => Cmult[18]) = "";
		(Bmult[8]  => Cmult[18]) = "";
		(Bmult[9]  => Cmult[18]) = "";
		(Bmult[10] => Cmult[18]) = "";
		(Bmult[11] => Cmult[18]) = "";
		(Bmult[12] => Cmult[18]) = "";
		(Bmult[13] => Cmult[18]) = "";
		(Bmult[14] => Cmult[18]) = "";
		(Bmult[15] => Cmult[18]) = "";
		(Bmult[16] => Cmult[18]) = "";
		(Bmult[17] => Cmult[18]) = "";
		(Bmult[18] => Cmult[18]) = "";
		(Bmult[19] => Cmult[18]) = "";
		(Bmult[20] => Cmult[18]) = "";
		(Bmult[21] => Cmult[18]) = "";
		(Bmult[22] => Cmult[18]) = "";
		(Bmult[23] => Cmult[18]) = "";
		(Bmult[24] => Cmult[18]) = "";
		(Bmult[25] => Cmult[18]) = "";
		(Bmult[26] => Cmult[18]) = "";
		(Bmult[27] => Cmult[18]) = "";
		(Bmult[28] => Cmult[18]) = "";
		(Bmult[29] => Cmult[18]) = "";
		(Bmult[30] => Cmult[18]) = "";
		(Bmult[31] => Cmult[18]) = "";		
		(Valid_mult[0] => Cmult[18]) = "";
		(Valid_mult[1] => Cmult[18]) = "";
		(sel_mul_32x32 => Cmult[18]) = "";	
		(Amult[0]  => Cmult[19]) = "";
		(Amult[1]  => Cmult[19]) = "";
		(Amult[2]  => Cmult[19]) = "";
		(Amult[3]  => Cmult[19]) = "";
		(Amult[4]  => Cmult[19]) = "";
		(Amult[5]  => Cmult[19]) = "";
		(Amult[6]  => Cmult[19]) = "";
		(Amult[7]  => Cmult[19]) = "";
		(Amult[8]  => Cmult[19]) = "";
		(Amult[9]  => Cmult[19]) = "";
		(Amult[10] => Cmult[19]) = "";
		(Amult[11] => Cmult[19]) = "";
		(Amult[12] => Cmult[19]) = "";
		(Amult[13] => Cmult[19]) = "";
		(Amult[14] => Cmult[19]) = "";
		(Amult[15] => Cmult[19]) = "";
		(Amult[16] => Cmult[19]) = "";
		(Amult[17] => Cmult[19]) = "";
		(Amult[18] => Cmult[19]) = "";
		(Amult[19] => Cmult[19]) = "";
		(Amult[20] => Cmult[19]) = "";
		(Amult[21] => Cmult[19]) = "";
		(Amult[22] => Cmult[19]) = "";
		(Amult[23] => Cmult[19]) = "";
		(Amult[24] => Cmult[19]) = "";
		(Amult[25] => Cmult[19]) = "";
		(Amult[26] => Cmult[19]) = "";
		(Amult[27] => Cmult[19]) = "";
		(Amult[28] => Cmult[19]) = "";
		(Amult[29] => Cmult[19]) = "";
		(Amult[30] => Cmult[19]) = "";
		(Amult[31] => Cmult[19]) = "";
		(Bmult[0]  => Cmult[19]) = "";
		(Bmult[1]  => Cmult[19]) = "";
		(Bmult[2]  => Cmult[19]) = "";
		(Bmult[3]  => Cmult[19]) = "";
		(Bmult[4]  => Cmult[19]) = "";
		(Bmult[5]  => Cmult[19]) = "";
		(Bmult[6]  => Cmult[19]) = "";
		(Bmult[7]  => Cmult[19]) = "";
		(Bmult[8]  => Cmult[19]) = "";
		(Bmult[9]  => Cmult[19]) = "";
		(Bmult[10] => Cmult[19]) = "";
		(Bmult[11] => Cmult[19]) = "";
		(Bmult[12] => Cmult[19]) = "";
		(Bmult[13] => Cmult[19]) = "";
		(Bmult[14] => Cmult[19]) = "";
		(Bmult[15] => Cmult[19]) = "";
		(Bmult[16] => Cmult[19]) = "";
		(Bmult[17] => Cmult[19]) = "";
		(Bmult[18] => Cmult[19]) = "";
		(Bmult[19] => Cmult[19]) = "";
		(Bmult[20] => Cmult[19]) = "";
		(Bmult[21] => Cmult[19]) = "";
		(Bmult[22] => Cmult[19]) = "";
		(Bmult[23] => Cmult[19]) = "";
		(Bmult[24] => Cmult[19]) = "";
		(Bmult[25] => Cmult[19]) = "";
		(Bmult[26] => Cmult[19]) = "";
		(Bmult[27] => Cmult[19]) = "";
		(Bmult[28] => Cmult[19]) = "";
		(Bmult[29] => Cmult[19]) = "";
		(Bmult[30] => Cmult[19]) = "";
		(Bmult[31] => Cmult[19]) = "";		
		(Valid_mult[0] => Cmult[19]) = "";
		(Valid_mult[1] => Cmult[19]) = "";
		(sel_mul_32x32 => Cmult[19]) = "";
		(Amult[0]  => Cmult[20]) = "";
		(Amult[1]  => Cmult[20]) = "";
		(Amult[2]  => Cmult[20]) = "";
		(Amult[3]  => Cmult[20]) = "";
		(Amult[4]  => Cmult[20]) = "";
		(Amult[5]  => Cmult[20]) = "";
		(Amult[6]  => Cmult[20]) = "";
		(Amult[7]  => Cmult[20]) = "";
		(Amult[8]  => Cmult[20]) = "";
		(Amult[9]  => Cmult[20]) = "";
		(Amult[10] => Cmult[20]) = "";
		(Amult[11] => Cmult[20]) = "";
		(Amult[12] => Cmult[20]) = "";
		(Amult[13] => Cmult[20]) = "";
		(Amult[14] => Cmult[20]) = "";
		(Amult[15] => Cmult[20]) = "";
		(Amult[16] => Cmult[20]) = "";
		(Amult[17] => Cmult[20]) = "";
		(Amult[18] => Cmult[20]) = "";
		(Amult[19] => Cmult[20]) = "";
		(Amult[20] => Cmult[20]) = "";
		(Amult[21] => Cmult[20]) = "";
		(Amult[22] => Cmult[20]) = "";
		(Amult[23] => Cmult[20]) = "";
		(Amult[24] => Cmult[20]) = "";
		(Amult[25] => Cmult[20]) = "";
		(Amult[26] => Cmult[20]) = "";
		(Amult[27] => Cmult[20]) = "";
		(Amult[28] => Cmult[20]) = "";
		(Amult[29] => Cmult[20]) = "";
		(Amult[30] => Cmult[20]) = "";
		(Amult[31] => Cmult[20]) = "";
		(Bmult[0]  => Cmult[20]) = "";
		(Bmult[1]  => Cmult[20]) = "";
		(Bmult[2]  => Cmult[20]) = "";
		(Bmult[3]  => Cmult[20]) = "";
		(Bmult[4]  => Cmult[20]) = "";
		(Bmult[5]  => Cmult[20]) = "";
		(Bmult[6]  => Cmult[20]) = "";
		(Bmult[7]  => Cmult[20]) = "";
		(Bmult[8]  => Cmult[20]) = "";
		(Bmult[9]  => Cmult[20]) = "";
		(Bmult[10] => Cmult[20]) = "";
		(Bmult[11] => Cmult[20]) = "";
		(Bmult[12] => Cmult[20]) = "";
		(Bmult[13] => Cmult[20]) = "";
		(Bmult[14] => Cmult[20]) = "";
		(Bmult[15] => Cmult[20]) = "";
		(Bmult[16] => Cmult[20]) = "";
		(Bmult[17] => Cmult[20]) = "";
		(Bmult[18] => Cmult[20]) = "";
		(Bmult[19] => Cmult[20]) = "";
		(Bmult[20] => Cmult[20]) = "";
		(Bmult[21] => Cmult[20]) = "";
		(Bmult[22] => Cmult[20]) = "";
		(Bmult[23] => Cmult[20]) = "";
		(Bmult[24] => Cmult[20]) = "";
		(Bmult[25] => Cmult[20]) = "";
		(Bmult[26] => Cmult[20]) = "";
		(Bmult[27] => Cmult[20]) = "";
		(Bmult[28] => Cmult[20]) = "";
		(Bmult[29] => Cmult[20]) = "";
		(Bmult[30] => Cmult[20]) = "";
		(Bmult[31] => Cmult[20]) = "";		
		(Valid_mult[0] => Cmult[20]) = "";
		(Valid_mult[1] => Cmult[20]) = "";
		(sel_mul_32x32 => Cmult[20]) = "";
		(Amult[0]  => Cmult[21]) = "";
		(Amult[1]  => Cmult[21]) = "";
		(Amult[2]  => Cmult[21]) = "";
		(Amult[3]  => Cmult[21]) = "";
		(Amult[4]  => Cmult[21]) = "";
		(Amult[5]  => Cmult[21]) = "";
		(Amult[6]  => Cmult[21]) = "";
		(Amult[7]  => Cmult[21]) = "";
		(Amult[8]  => Cmult[21]) = "";
		(Amult[9]  => Cmult[21]) = "";
		(Amult[10] => Cmult[21]) = "";
		(Amult[11] => Cmult[21]) = "";
		(Amult[12] => Cmult[21]) = "";
		(Amult[13] => Cmult[21]) = "";
		(Amult[14] => Cmult[21]) = "";
		(Amult[15] => Cmult[21]) = "";
		(Amult[16] => Cmult[21]) = "";
		(Amult[17] => Cmult[21]) = "";
		(Amult[18] => Cmult[21]) = "";
		(Amult[19] => Cmult[21]) = "";
		(Amult[20] => Cmult[21]) = "";
		(Amult[21] => Cmult[21]) = "";
		(Amult[22] => Cmult[21]) = "";
		(Amult[23] => Cmult[21]) = "";
		(Amult[24] => Cmult[21]) = "";
		(Amult[25] => Cmult[21]) = "";
		(Amult[26] => Cmult[21]) = "";
		(Amult[27] => Cmult[21]) = "";
		(Amult[28] => Cmult[21]) = "";
		(Amult[29] => Cmult[21]) = "";
		(Amult[30] => Cmult[21]) = "";
		(Amult[31] => Cmult[21]) = "";
		(Bmult[0]  => Cmult[21]) = "";
		(Bmult[1]  => Cmult[21]) = "";
		(Bmult[2]  => Cmult[21]) = "";
		(Bmult[3]  => Cmult[21]) = "";
		(Bmult[4]  => Cmult[21]) = "";
		(Bmult[5]  => Cmult[21]) = "";
		(Bmult[6]  => Cmult[21]) = "";
		(Bmult[7]  => Cmult[21]) = "";
		(Bmult[8]  => Cmult[21]) = "";
		(Bmult[9]  => Cmult[21]) = "";
		(Bmult[10] => Cmult[21]) = "";
		(Bmult[11] => Cmult[21]) = "";
		(Bmult[12] => Cmult[21]) = "";
		(Bmult[13] => Cmult[21]) = "";
		(Bmult[14] => Cmult[21]) = "";
		(Bmult[15] => Cmult[21]) = "";
		(Bmult[16] => Cmult[21]) = "";
		(Bmult[17] => Cmult[21]) = "";
		(Bmult[18] => Cmult[21]) = "";
		(Bmult[19] => Cmult[21]) = "";
		(Bmult[20] => Cmult[21]) = "";
		(Bmult[21] => Cmult[21]) = "";
		(Bmult[22] => Cmult[21]) = "";
		(Bmult[23] => Cmult[21]) = "";
		(Bmult[24] => Cmult[21]) = "";
		(Bmult[25] => Cmult[21]) = "";
		(Bmult[26] => Cmult[21]) = "";
		(Bmult[27] => Cmult[21]) = "";
		(Bmult[28] => Cmult[21]) = "";
		(Bmult[29] => Cmult[21]) = "";
		(Bmult[30] => Cmult[21]) = "";
		(Bmult[31] => Cmult[21]) = "";		
		(Valid_mult[0] => Cmult[21]) = "";
		(Valid_mult[1] => Cmult[21]) = "";
		(sel_mul_32x32 => Cmult[21]) = "";
		(Amult[0]  => Cmult[22]) = "";
		(Amult[1]  => Cmult[22]) = "";
		(Amult[2]  => Cmult[22]) = "";
		(Amult[3]  => Cmult[22]) = "";
		(Amult[4]  => Cmult[22]) = "";
		(Amult[5]  => Cmult[22]) = "";
		(Amult[6]  => Cmult[22]) = "";
		(Amult[7]  => Cmult[22]) = "";
		(Amult[8]  => Cmult[22]) = "";
		(Amult[9]  => Cmult[22]) = "";
		(Amult[10] => Cmult[22]) = "";
		(Amult[11] => Cmult[22]) = "";
		(Amult[12] => Cmult[22]) = "";
		(Amult[13] => Cmult[22]) = "";
		(Amult[14] => Cmult[22]) = "";
		(Amult[15] => Cmult[22]) = "";
		(Amult[16] => Cmult[22]) = "";
		(Amult[17] => Cmult[22]) = "";
		(Amult[18] => Cmult[22]) = "";
		(Amult[19] => Cmult[22]) = "";
		(Amult[20] => Cmult[22]) = "";
		(Amult[21] => Cmult[22]) = "";
		(Amult[22] => Cmult[22]) = "";
		(Amult[23] => Cmult[22]) = "";
		(Amult[24] => Cmult[22]) = "";
		(Amult[25] => Cmult[22]) = "";
		(Amult[26] => Cmult[22]) = "";
		(Amult[27] => Cmult[22]) = "";
		(Amult[28] => Cmult[22]) = "";
		(Amult[29] => Cmult[22]) = "";
		(Amult[30] => Cmult[22]) = "";
		(Amult[31] => Cmult[22]) = "";
		(Bmult[0]  => Cmult[22]) = "";
		(Bmult[1]  => Cmult[22]) = "";
		(Bmult[2]  => Cmult[22]) = "";
		(Bmult[3]  => Cmult[22]) = "";
		(Bmult[4]  => Cmult[22]) = "";
		(Bmult[5]  => Cmult[22]) = "";
		(Bmult[6]  => Cmult[22]) = "";
		(Bmult[7]  => Cmult[22]) = "";
		(Bmult[8]  => Cmult[22]) = "";
		(Bmult[9]  => Cmult[22]) = "";
		(Bmult[10] => Cmult[22]) = "";
		(Bmult[11] => Cmult[22]) = "";
		(Bmult[12] => Cmult[22]) = "";
		(Bmult[13] => Cmult[22]) = "";
		(Bmult[14] => Cmult[22]) = "";
		(Bmult[15] => Cmult[22]) = "";
		(Bmult[16] => Cmult[22]) = "";
		(Bmult[17] => Cmult[22]) = "";
		(Bmult[18] => Cmult[22]) = "";
		(Bmult[19] => Cmult[22]) = "";
		(Bmult[20] => Cmult[22]) = "";
		(Bmult[21] => Cmult[22]) = "";
		(Bmult[22] => Cmult[22]) = "";
		(Bmult[23] => Cmult[22]) = "";
		(Bmult[24] => Cmult[22]) = "";
		(Bmult[25] => Cmult[22]) = "";
		(Bmult[26] => Cmult[22]) = "";
		(Bmult[27] => Cmult[22]) = "";
		(Bmult[28] => Cmult[22]) = "";
		(Bmult[29] => Cmult[22]) = "";
		(Bmult[30] => Cmult[22]) = "";
		(Bmult[31] => Cmult[22]) = "";		
		(Valid_mult[0] => Cmult[22]) = "";
		(Valid_mult[1] => Cmult[22]) = "";
		(sel_mul_32x32 => Cmult[22]) = "";
		(Amult[0]  => Cmult[23]) = "";
		(Amult[1]  => Cmult[23]) = "";
		(Amult[2]  => Cmult[23]) = "";
		(Amult[3]  => Cmult[23]) = "";
		(Amult[4]  => Cmult[23]) = "";
		(Amult[5]  => Cmult[23]) = "";
		(Amult[6]  => Cmult[23]) = "";
		(Amult[7]  => Cmult[23]) = "";
		(Amult[8]  => Cmult[23]) = "";
		(Amult[9]  => Cmult[23]) = "";
		(Amult[10] => Cmult[23]) = "";
		(Amult[11] => Cmult[23]) = "";
		(Amult[12] => Cmult[23]) = "";
		(Amult[13] => Cmult[23]) = "";
		(Amult[14] => Cmult[23]) = "";
		(Amult[15] => Cmult[23]) = "";
		(Amult[16] => Cmult[23]) = "";
		(Amult[17] => Cmult[23]) = "";
		(Amult[18] => Cmult[23]) = "";
		(Amult[19] => Cmult[23]) = "";
		(Amult[20] => Cmult[23]) = "";
		(Amult[21] => Cmult[23]) = "";
		(Amult[22] => Cmult[23]) = "";
		(Amult[23] => Cmult[23]) = "";
		(Amult[24] => Cmult[23]) = "";
		(Amult[25] => Cmult[23]) = "";
		(Amult[26] => Cmult[23]) = "";
		(Amult[27] => Cmult[23]) = "";
		(Amult[28] => Cmult[23]) = "";
		(Amult[29] => Cmult[23]) = "";
		(Amult[30] => Cmult[23]) = "";
		(Amult[31] => Cmult[23]) = "";
		(Bmult[0]  => Cmult[23]) = "";
		(Bmult[1]  => Cmult[23]) = "";
		(Bmult[2]  => Cmult[23]) = "";
		(Bmult[3]  => Cmult[23]) = "";
		(Bmult[4]  => Cmult[23]) = "";
		(Bmult[5]  => Cmult[23]) = "";
		(Bmult[6]  => Cmult[23]) = "";
		(Bmult[7]  => Cmult[23]) = "";
		(Bmult[8]  => Cmult[23]) = "";
		(Bmult[9]  => Cmult[23]) = "";
		(Bmult[10] => Cmult[23]) = "";
		(Bmult[11] => Cmult[23]) = "";
		(Bmult[12] => Cmult[23]) = "";
		(Bmult[13] => Cmult[23]) = "";
		(Bmult[14] => Cmult[23]) = "";
		(Bmult[15] => Cmult[23]) = "";
		(Bmult[16] => Cmult[23]) = "";
		(Bmult[17] => Cmult[23]) = "";
		(Bmult[18] => Cmult[23]) = "";
		(Bmult[19] => Cmult[23]) = "";
		(Bmult[20] => Cmult[23]) = "";
		(Bmult[21] => Cmult[23]) = "";
		(Bmult[22] => Cmult[23]) = "";
		(Bmult[23] => Cmult[23]) = "";
		(Bmult[24] => Cmult[23]) = "";
		(Bmult[25] => Cmult[23]) = "";
		(Bmult[26] => Cmult[23]) = "";
		(Bmult[27] => Cmult[23]) = "";
		(Bmult[28] => Cmult[23]) = "";
		(Bmult[29] => Cmult[23]) = "";
		(Bmult[30] => Cmult[23]) = "";
		(Bmult[31] => Cmult[23]) = "";		
		(Valid_mult[0] => Cmult[23]) = "";
		(Valid_mult[1] => Cmult[23]) = "";
		(sel_mul_32x32 => Cmult[23]) = "";
		(Amult[0]  => Cmult[24]) = "";
		(Amult[1]  => Cmult[24]) = "";
		(Amult[2]  => Cmult[24]) = "";
		(Amult[3]  => Cmult[24]) = "";
		(Amult[4]  => Cmult[24]) = "";
		(Amult[5]  => Cmult[24]) = "";
		(Amult[6]  => Cmult[24]) = "";
		(Amult[7]  => Cmult[24]) = "";
		(Amult[8]  => Cmult[24]) = "";
		(Amult[9]  => Cmult[24]) = "";
		(Amult[10] => Cmult[24]) = "";
		(Amult[11] => Cmult[24]) = "";
		(Amult[12] => Cmult[24]) = "";
		(Amult[13] => Cmult[24]) = "";
		(Amult[14] => Cmult[24]) = "";
		(Amult[15] => Cmult[24]) = "";
		(Amult[16] => Cmult[24]) = "";
		(Amult[17] => Cmult[24]) = "";
		(Amult[18] => Cmult[24]) = "";
		(Amult[19] => Cmult[24]) = "";
		(Amult[20] => Cmult[24]) = "";
		(Amult[21] => Cmult[24]) = "";
		(Amult[22] => Cmult[24]) = "";
		(Amult[23] => Cmult[24]) = "";
		(Amult[24] => Cmult[24]) = "";
		(Amult[25] => Cmult[24]) = "";
		(Amult[26] => Cmult[24]) = "";
		(Amult[27] => Cmult[24]) = "";
		(Amult[28] => Cmult[24]) = "";
		(Amult[29] => Cmult[24]) = "";
		(Amult[30] => Cmult[24]) = "";
		(Amult[31] => Cmult[24]) = "";
		(Bmult[0]  => Cmult[24]) = "";
		(Bmult[1]  => Cmult[24]) = "";
		(Bmult[2]  => Cmult[24]) = "";
		(Bmult[3]  => Cmult[24]) = "";
		(Bmult[4]  => Cmult[24]) = "";
		(Bmult[5]  => Cmult[24]) = "";
		(Bmult[6]  => Cmult[24]) = "";
		(Bmult[7]  => Cmult[24]) = "";
		(Bmult[8]  => Cmult[24]) = "";
		(Bmult[9]  => Cmult[24]) = "";
		(Bmult[10] => Cmult[24]) = "";
		(Bmult[11] => Cmult[24]) = "";
		(Bmult[12] => Cmult[24]) = "";
		(Bmult[13] => Cmult[24]) = "";
		(Bmult[14] => Cmult[24]) = "";
		(Bmult[15] => Cmult[24]) = "";
		(Bmult[16] => Cmult[24]) = "";
		(Bmult[17] => Cmult[24]) = "";
		(Bmult[18] => Cmult[24]) = "";
		(Bmult[19] => Cmult[24]) = "";
		(Bmult[20] => Cmult[24]) = "";
		(Bmult[21] => Cmult[24]) = "";
		(Bmult[22] => Cmult[24]) = "";
		(Bmult[23] => Cmult[24]) = "";
		(Bmult[24] => Cmult[24]) = "";
		(Bmult[25] => Cmult[24]) = "";
		(Bmult[26] => Cmult[24]) = "";
		(Bmult[27] => Cmult[24]) = "";
		(Bmult[28] => Cmult[24]) = "";
		(Bmult[29] => Cmult[24]) = "";
		(Bmult[30] => Cmult[24]) = "";
		(Bmult[31] => Cmult[24]) = "";		
		(Valid_mult[0] => Cmult[24]) = "";
		(Valid_mult[1] => Cmult[24]) = "";
		(sel_mul_32x32 => Cmult[24]) = "";
		(Amult[0]  => Cmult[25]) = "";
		(Amult[1]  => Cmult[25]) = "";
		(Amult[2]  => Cmult[25]) = "";
		(Amult[3]  => Cmult[25]) = "";
		(Amult[4]  => Cmult[25]) = "";
		(Amult[5]  => Cmult[25]) = "";
		(Amult[6]  => Cmult[25]) = "";
		(Amult[7]  => Cmult[25]) = "";
		(Amult[8]  => Cmult[25]) = "";
		(Amult[9]  => Cmult[25]) = "";
		(Amult[10] => Cmult[25]) = "";
		(Amult[11] => Cmult[25]) = "";
		(Amult[12] => Cmult[25]) = "";
		(Amult[13] => Cmult[25]) = "";
		(Amult[14] => Cmult[25]) = "";
		(Amult[15] => Cmult[25]) = "";
		(Amult[16] => Cmult[25]) = "";
		(Amult[17] => Cmult[25]) = "";
		(Amult[18] => Cmult[25]) = "";
		(Amult[19] => Cmult[25]) = "";
		(Amult[20] => Cmult[25]) = "";
		(Amult[21] => Cmult[25]) = "";
		(Amult[22] => Cmult[25]) = "";
		(Amult[23] => Cmult[25]) = "";
		(Amult[24] => Cmult[25]) = "";
		(Amult[25] => Cmult[25]) = "";
		(Amult[26] => Cmult[25]) = "";
		(Amult[27] => Cmult[25]) = "";
		(Amult[28] => Cmult[25]) = "";
		(Amult[29] => Cmult[25]) = "";
		(Amult[30] => Cmult[25]) = "";
		(Amult[31] => Cmult[25]) = "";
		(Bmult[0]  => Cmult[25]) = "";
		(Bmult[1]  => Cmult[25]) = "";
		(Bmult[2]  => Cmult[25]) = "";
		(Bmult[3]  => Cmult[25]) = "";
		(Bmult[4]  => Cmult[25]) = "";
		(Bmult[5]  => Cmult[25]) = "";
		(Bmult[6]  => Cmult[25]) = "";
		(Bmult[7]  => Cmult[25]) = "";
		(Bmult[8]  => Cmult[25]) = "";
		(Bmult[9]  => Cmult[25]) = "";
		(Bmult[10] => Cmult[25]) = "";
		(Bmult[11] => Cmult[25]) = "";
		(Bmult[12] => Cmult[25]) = "";
		(Bmult[13] => Cmult[25]) = "";
		(Bmult[14] => Cmult[25]) = "";
		(Bmult[15] => Cmult[25]) = "";
		(Bmult[16] => Cmult[25]) = "";
		(Bmult[17] => Cmult[25]) = "";
		(Bmult[18] => Cmult[25]) = "";
		(Bmult[19] => Cmult[25]) = "";
		(Bmult[20] => Cmult[25]) = "";
		(Bmult[21] => Cmult[25]) = "";
		(Bmult[22] => Cmult[25]) = "";
		(Bmult[23] => Cmult[25]) = "";
		(Bmult[24] => Cmult[25]) = "";
		(Bmult[25] => Cmult[25]) = "";
		(Bmult[26] => Cmult[25]) = "";
		(Bmult[27] => Cmult[25]) = "";
		(Bmult[28] => Cmult[25]) = "";
		(Bmult[29] => Cmult[25]) = "";
		(Bmult[30] => Cmult[25]) = "";
		(Bmult[31] => Cmult[25]) = "";		
		(Valid_mult[0] => Cmult[25]) = "";
		(Valid_mult[1] => Cmult[25]) = "";
		(sel_mul_32x32 => Cmult[25]) = "";
		(Amult[0]  => Cmult[26]) = "";
		(Amult[1]  => Cmult[26]) = "";
		(Amult[2]  => Cmult[26]) = "";
		(Amult[3]  => Cmult[26]) = "";
		(Amult[4]  => Cmult[26]) = "";
		(Amult[5]  => Cmult[26]) = "";
		(Amult[6]  => Cmult[26]) = "";
		(Amult[7]  => Cmult[26]) = "";
		(Amult[8]  => Cmult[26]) = "";
		(Amult[9]  => Cmult[26]) = "";
		(Amult[10] => Cmult[26]) = "";
		(Amult[11] => Cmult[26]) = "";
		(Amult[12] => Cmult[26]) = "";
		(Amult[13] => Cmult[26]) = "";
		(Amult[14] => Cmult[26]) = "";
		(Amult[15] => Cmult[26]) = "";
		(Amult[16] => Cmult[26]) = "";
		(Amult[17] => Cmult[26]) = "";
		(Amult[18] => Cmult[26]) = "";
		(Amult[19] => Cmult[26]) = "";
		(Amult[20] => Cmult[26]) = "";
		(Amult[21] => Cmult[26]) = "";
		(Amult[22] => Cmult[26]) = "";
		(Amult[23] => Cmult[26]) = "";
		(Amult[24] => Cmult[26]) = "";
		(Amult[25] => Cmult[26]) = "";
		(Amult[26] => Cmult[26]) = "";
		(Amult[27] => Cmult[26]) = "";
		(Amult[28] => Cmult[26]) = "";
		(Amult[29] => Cmult[26]) = "";
		(Amult[30] => Cmult[26]) = "";
		(Amult[31] => Cmult[26]) = "";
		(Bmult[0]  => Cmult[26]) = "";
		(Bmult[1]  => Cmult[26]) = "";
		(Bmult[2]  => Cmult[26]) = "";
		(Bmult[3]  => Cmult[26]) = "";
		(Bmult[4]  => Cmult[26]) = "";
		(Bmult[5]  => Cmult[26]) = "";
		(Bmult[6]  => Cmult[26]) = "";
		(Bmult[7]  => Cmult[26]) = "";
		(Bmult[8]  => Cmult[26]) = "";
		(Bmult[9]  => Cmult[26]) = "";
		(Bmult[10] => Cmult[26]) = "";
		(Bmult[11] => Cmult[26]) = "";
		(Bmult[12] => Cmult[26]) = "";
		(Bmult[13] => Cmult[26]) = "";
		(Bmult[14] => Cmult[26]) = "";
		(Bmult[15] => Cmult[26]) = "";
		(Bmult[16] => Cmult[26]) = "";
		(Bmult[17] => Cmult[26]) = "";
		(Bmult[18] => Cmult[26]) = "";
		(Bmult[19] => Cmult[26]) = "";
		(Bmult[20] => Cmult[26]) = "";
		(Bmult[21] => Cmult[26]) = "";
		(Bmult[22] => Cmult[26]) = "";
		(Bmult[23] => Cmult[26]) = "";
		(Bmult[24] => Cmult[26]) = "";
		(Bmult[25] => Cmult[26]) = "";
		(Bmult[26] => Cmult[26]) = "";
		(Bmult[27] => Cmult[26]) = "";
		(Bmult[28] => Cmult[26]) = "";
		(Bmult[29] => Cmult[26]) = "";
		(Bmult[30] => Cmult[26]) = "";
		(Bmult[31] => Cmult[26]) = "";		
		(Valid_mult[0] => Cmult[26]) = "";
		(Valid_mult[1] => Cmult[26]) = "";
		(sel_mul_32x32 => Cmult[26]) = "";
		(Amult[0]  => Cmult[27]) = "";
		(Amult[1]  => Cmult[27]) = "";
		(Amult[2]  => Cmult[27]) = "";
		(Amult[3]  => Cmult[27]) = "";
		(Amult[4]  => Cmult[27]) = "";
		(Amult[5]  => Cmult[27]) = "";
		(Amult[6]  => Cmult[27]) = "";
		(Amult[7]  => Cmult[27]) = "";
		(Amult[8]  => Cmult[27]) = "";
		(Amult[9]  => Cmult[27]) = "";
		(Amult[10] => Cmult[27]) = "";
		(Amult[11] => Cmult[27]) = "";
		(Amult[12] => Cmult[27]) = "";
		(Amult[13] => Cmult[27]) = "";
		(Amult[14] => Cmult[27]) = "";
		(Amult[15] => Cmult[27]) = "";
		(Amult[16] => Cmult[27]) = "";
		(Amult[17] => Cmult[27]) = "";
		(Amult[18] => Cmult[27]) = "";
		(Amult[19] => Cmult[27]) = "";
		(Amult[20] => Cmult[27]) = "";
		(Amult[21] => Cmult[27]) = "";
		(Amult[22] => Cmult[27]) = "";
		(Amult[23] => Cmult[27]) = "";
		(Amult[24] => Cmult[27]) = "";
		(Amult[25] => Cmult[27]) = "";
		(Amult[26] => Cmult[27]) = "";
		(Amult[27] => Cmult[27]) = "";
		(Amult[28] => Cmult[27]) = "";
		(Amult[29] => Cmult[27]) = "";
		(Amult[30] => Cmult[27]) = "";
		(Amult[31] => Cmult[27]) = "";
		(Bmult[0]  => Cmult[27]) = "";
		(Bmult[1]  => Cmult[27]) = "";
		(Bmult[2]  => Cmult[27]) = "";
		(Bmult[3]  => Cmult[27]) = "";
		(Bmult[4]  => Cmult[27]) = "";
		(Bmult[5]  => Cmult[27]) = "";
		(Bmult[6]  => Cmult[27]) = "";
		(Bmult[7]  => Cmult[27]) = "";
		(Bmult[8]  => Cmult[27]) = "";
		(Bmult[9]  => Cmult[27]) = "";
		(Bmult[10] => Cmult[27]) = "";
		(Bmult[11] => Cmult[27]) = "";
		(Bmult[12] => Cmult[27]) = "";
		(Bmult[13] => Cmult[27]) = "";
		(Bmult[14] => Cmult[27]) = "";
		(Bmult[15] => Cmult[27]) = "";
		(Bmult[16] => Cmult[27]) = "";
		(Bmult[17] => Cmult[27]) = "";
		(Bmult[18] => Cmult[27]) = "";
		(Bmult[19] => Cmult[27]) = "";
		(Bmult[20] => Cmult[27]) = "";
		(Bmult[21] => Cmult[27]) = "";
		(Bmult[22] => Cmult[27]) = "";
		(Bmult[23] => Cmult[27]) = "";
		(Bmult[24] => Cmult[27]) = "";
		(Bmult[25] => Cmult[27]) = "";
		(Bmult[26] => Cmult[27]) = "";
		(Bmult[27] => Cmult[27]) = "";
		(Bmult[28] => Cmult[27]) = "";
		(Bmult[29] => Cmult[27]) = "";
		(Bmult[30] => Cmult[27]) = "";
		(Bmult[31] => Cmult[27]) = "";		
		(Valid_mult[0] => Cmult[27]) = "";
		(Valid_mult[1] => Cmult[27]) = "";
		(sel_mul_32x32 => Cmult[27]) = "";
		(Amult[0]  => Cmult[28]) = "";
		(Amult[1]  => Cmult[28]) = "";
		(Amult[2]  => Cmult[28]) = "";
		(Amult[3]  => Cmult[28]) = "";
		(Amult[4]  => Cmult[28]) = "";
		(Amult[5]  => Cmult[28]) = "";
		(Amult[6]  => Cmult[28]) = "";
		(Amult[7]  => Cmult[28]) = "";
		(Amult[8]  => Cmult[28]) = "";
		(Amult[9]  => Cmult[28]) = "";
		(Amult[10] => Cmult[28]) = "";
		(Amult[11] => Cmult[28]) = "";
		(Amult[12] => Cmult[28]) = "";
		(Amult[13] => Cmult[28]) = "";
		(Amult[14] => Cmult[28]) = "";
		(Amult[15] => Cmult[28]) = "";
		(Amult[16] => Cmult[28]) = "";
		(Amult[17] => Cmult[28]) = "";
		(Amult[18] => Cmult[28]) = "";
		(Amult[19] => Cmult[28]) = "";
		(Amult[20] => Cmult[28]) = "";
		(Amult[21] => Cmult[28]) = "";
		(Amult[22] => Cmult[28]) = "";
		(Amult[23] => Cmult[28]) = "";
		(Amult[24] => Cmult[28]) = "";
		(Amult[25] => Cmult[28]) = "";
		(Amult[26] => Cmult[28]) = "";
		(Amult[27] => Cmult[28]) = "";
		(Amult[28] => Cmult[28]) = "";
		(Amult[29] => Cmult[28]) = "";
		(Amult[30] => Cmult[28]) = "";
		(Amult[31] => Cmult[28]) = "";
		(Bmult[0]  => Cmult[28]) = "";
		(Bmult[1]  => Cmult[28]) = "";
		(Bmult[2]  => Cmult[28]) = "";
		(Bmult[3]  => Cmult[28]) = "";
		(Bmult[4]  => Cmult[28]) = "";
		(Bmult[5]  => Cmult[28]) = "";
		(Bmult[6]  => Cmult[28]) = "";
		(Bmult[7]  => Cmult[28]) = "";
		(Bmult[8]  => Cmult[28]) = "";
		(Bmult[9]  => Cmult[28]) = "";
		(Bmult[10] => Cmult[28]) = "";
		(Bmult[11] => Cmult[28]) = "";
		(Bmult[12] => Cmult[28]) = "";
		(Bmult[13] => Cmult[28]) = "";
		(Bmult[14] => Cmult[28]) = "";
		(Bmult[15] => Cmult[28]) = "";
		(Bmult[16] => Cmult[28]) = "";
		(Bmult[17] => Cmult[28]) = "";
		(Bmult[18] => Cmult[28]) = "";
		(Bmult[19] => Cmult[28]) = "";
		(Bmult[20] => Cmult[28]) = "";
		(Bmult[21] => Cmult[28]) = "";
		(Bmult[22] => Cmult[28]) = "";
		(Bmult[23] => Cmult[28]) = "";
		(Bmult[24] => Cmult[28]) = "";
		(Bmult[25] => Cmult[28]) = "";
		(Bmult[26] => Cmult[28]) = "";
		(Bmult[27] => Cmult[28]) = "";
		(Bmult[28] => Cmult[28]) = "";
		(Bmult[29] => Cmult[28]) = "";
		(Bmult[30] => Cmult[28]) = "";
		(Bmult[31] => Cmult[28]) = "";		
		(Valid_mult[0] => Cmult[28]) = "";
		(Valid_mult[1] => Cmult[28]) = "";
		(sel_mul_32x32 => Cmult[28]) = "";	
		(Amult[0]  => Cmult[29]) = "";
		(Amult[1]  => Cmult[29]) = "";
		(Amult[2]  => Cmult[29]) = "";
		(Amult[3]  => Cmult[29]) = "";
		(Amult[4]  => Cmult[29]) = "";
		(Amult[5]  => Cmult[29]) = "";
		(Amult[6]  => Cmult[29]) = "";
		(Amult[7]  => Cmult[29]) = "";
		(Amult[8]  => Cmult[29]) = "";
		(Amult[9]  => Cmult[29]) = "";
		(Amult[10] => Cmult[29]) = "";
		(Amult[11] => Cmult[29]) = "";
		(Amult[12] => Cmult[29]) = "";
		(Amult[13] => Cmult[29]) = "";
		(Amult[14] => Cmult[29]) = "";
		(Amult[15] => Cmult[29]) = "";
		(Amult[16] => Cmult[29]) = "";
		(Amult[17] => Cmult[29]) = "";
		(Amult[18] => Cmult[29]) = "";
		(Amult[19] => Cmult[29]) = "";
		(Amult[20] => Cmult[29]) = "";
		(Amult[21] => Cmult[29]) = "";
		(Amult[22] => Cmult[29]) = "";
		(Amult[23] => Cmult[29]) = "";
		(Amult[24] => Cmult[29]) = "";
		(Amult[25] => Cmult[29]) = "";
		(Amult[26] => Cmult[29]) = "";
		(Amult[27] => Cmult[29]) = "";
		(Amult[28] => Cmult[29]) = "";
		(Amult[29] => Cmult[29]) = "";
		(Amult[30] => Cmult[29]) = "";
		(Amult[31] => Cmult[29]) = "";
		(Bmult[0]  => Cmult[29]) = "";
		(Bmult[1]  => Cmult[29]) = "";
		(Bmult[2]  => Cmult[29]) = "";
		(Bmult[3]  => Cmult[29]) = "";
		(Bmult[4]  => Cmult[29]) = "";
		(Bmult[5]  => Cmult[29]) = "";
		(Bmult[6]  => Cmult[29]) = "";
		(Bmult[7]  => Cmult[29]) = "";
		(Bmult[8]  => Cmult[29]) = "";
		(Bmult[9]  => Cmult[29]) = "";
		(Bmult[10] => Cmult[29]) = "";
		(Bmult[11] => Cmult[29]) = "";
		(Bmult[12] => Cmult[29]) = "";
		(Bmult[13] => Cmult[29]) = "";
		(Bmult[14] => Cmult[29]) = "";
		(Bmult[15] => Cmult[29]) = "";
		(Bmult[16] => Cmult[29]) = "";
		(Bmult[17] => Cmult[29]) = "";
		(Bmult[18] => Cmult[29]) = "";
		(Bmult[19] => Cmult[29]) = "";
		(Bmult[20] => Cmult[29]) = "";
		(Bmult[21] => Cmult[29]) = "";
		(Bmult[22] => Cmult[29]) = "";
		(Bmult[23] => Cmult[29]) = "";
		(Bmult[24] => Cmult[29]) = "";
		(Bmult[25] => Cmult[29]) = "";
		(Bmult[26] => Cmult[29]) = "";
		(Bmult[27] => Cmult[29]) = "";
		(Bmult[28] => Cmult[29]) = "";
		(Bmult[29] => Cmult[29]) = "";
		(Bmult[30] => Cmult[29]) = "";
		(Bmult[31] => Cmult[29]) = "";		
		(Valid_mult[0] => Cmult[29]) = "";
		(Valid_mult[1] => Cmult[29]) = "";
		(sel_mul_32x32 => Cmult[29]) = "";	
		(Amult[0]  => Cmult[30]) = "";
		(Amult[1]  => Cmult[30]) = "";
		(Amult[2]  => Cmult[30]) = "";
		(Amult[3]  => Cmult[30]) = "";
		(Amult[4]  => Cmult[30]) = "";
		(Amult[5]  => Cmult[30]) = "";
		(Amult[6]  => Cmult[30]) = "";
		(Amult[7]  => Cmult[30]) = "";
		(Amult[8]  => Cmult[30]) = "";
		(Amult[9]  => Cmult[30]) = "";
		(Amult[10] => Cmult[30]) = "";
		(Amult[11] => Cmult[30]) = "";
		(Amult[12] => Cmult[30]) = "";
		(Amult[13] => Cmult[30]) = "";
		(Amult[14] => Cmult[30]) = "";
		(Amult[15] => Cmult[30]) = "";
		(Amult[16] => Cmult[30]) = "";
		(Amult[17] => Cmult[30]) = "";
		(Amult[18] => Cmult[30]) = "";
		(Amult[19] => Cmult[30]) = "";
		(Amult[20] => Cmult[30]) = "";
		(Amult[21] => Cmult[30]) = "";
		(Amult[22] => Cmult[30]) = "";
		(Amult[23] => Cmult[30]) = "";
		(Amult[24] => Cmult[30]) = "";
		(Amult[25] => Cmult[30]) = "";
		(Amult[26] => Cmult[30]) = "";
		(Amult[27] => Cmult[30]) = "";
		(Amult[28] => Cmult[30]) = "";
		(Amult[29] => Cmult[30]) = "";
		(Amult[30] => Cmult[30]) = "";
		(Amult[31] => Cmult[30]) = "";
		(Bmult[0]  => Cmult[30]) = "";
		(Bmult[1]  => Cmult[30]) = "";
		(Bmult[2]  => Cmult[30]) = "";
		(Bmult[3]  => Cmult[30]) = "";
		(Bmult[4]  => Cmult[30]) = "";
		(Bmult[5]  => Cmult[30]) = "";
		(Bmult[6]  => Cmult[30]) = "";
		(Bmult[7]  => Cmult[30]) = "";
		(Bmult[8]  => Cmult[30]) = "";
		(Bmult[9]  => Cmult[30]) = "";
		(Bmult[10] => Cmult[30]) = "";
		(Bmult[11] => Cmult[30]) = "";
		(Bmult[12] => Cmult[30]) = "";
		(Bmult[13] => Cmult[30]) = "";
		(Bmult[14] => Cmult[30]) = "";
		(Bmult[15] => Cmult[30]) = "";
		(Bmult[16] => Cmult[30]) = "";
		(Bmult[17] => Cmult[30]) = "";
		(Bmult[18] => Cmult[30]) = "";
		(Bmult[19] => Cmult[30]) = "";
		(Bmult[20] => Cmult[30]) = "";
		(Bmult[21] => Cmult[30]) = "";
		(Bmult[22] => Cmult[30]) = "";
		(Bmult[23] => Cmult[30]) = "";
		(Bmult[24] => Cmult[30]) = "";
		(Bmult[25] => Cmult[30]) = "";
		(Bmult[26] => Cmult[30]) = "";
		(Bmult[27] => Cmult[30]) = "";
		(Bmult[28] => Cmult[30]) = "";
		(Bmult[29] => Cmult[30]) = "";
		(Bmult[30] => Cmult[30]) = "";
		(Bmult[31] => Cmult[30]) = "";		
		(Valid_mult[0] => Cmult[30]) = "";
		(Valid_mult[1] => Cmult[30]) = "";
		(sel_mul_32x32 => Cmult[30]) = "";
		(Amult[0]  => Cmult[31]) = "";
		(Amult[1]  => Cmult[31]) = "";
		(Amult[2]  => Cmult[31]) = "";
		(Amult[3]  => Cmult[31]) = "";
		(Amult[4]  => Cmult[31]) = "";
		(Amult[5]  => Cmult[31]) = "";
		(Amult[6]  => Cmult[31]) = "";
		(Amult[7]  => Cmult[31]) = "";
		(Amult[8]  => Cmult[31]) = "";
		(Amult[9]  => Cmult[31]) = "";
		(Amult[10] => Cmult[31]) = "";
		(Amult[11] => Cmult[31]) = "";
		(Amult[12] => Cmult[31]) = "";
		(Amult[13] => Cmult[31]) = "";
		(Amult[14] => Cmult[31]) = "";
		(Amult[15] => Cmult[31]) = "";
		(Amult[16] => Cmult[31]) = "";
		(Amult[17] => Cmult[31]) = "";
		(Amult[18] => Cmult[31]) = "";
		(Amult[19] => Cmult[31]) = "";
		(Amult[20] => Cmult[31]) = "";
		(Amult[21] => Cmult[31]) = "";
		(Amult[22] => Cmult[31]) = "";
		(Amult[23] => Cmult[31]) = "";
		(Amult[24] => Cmult[31]) = "";
		(Amult[25] => Cmult[31]) = "";
		(Amult[26] => Cmult[31]) = "";
		(Amult[27] => Cmult[31]) = "";
		(Amult[28] => Cmult[31]) = "";
		(Amult[29] => Cmult[31]) = "";
		(Amult[30] => Cmult[31]) = "";
		(Amult[31] => Cmult[31]) = "";
		(Bmult[0]  => Cmult[31]) = "";
		(Bmult[1]  => Cmult[31]) = "";
		(Bmult[2]  => Cmult[31]) = "";
		(Bmult[3]  => Cmult[31]) = "";
		(Bmult[4]  => Cmult[31]) = "";
		(Bmult[5]  => Cmult[31]) = "";
		(Bmult[6]  => Cmult[31]) = "";
		(Bmult[7]  => Cmult[31]) = "";
		(Bmult[8]  => Cmult[31]) = "";
		(Bmult[9]  => Cmult[31]) = "";
		(Bmult[10] => Cmult[31]) = "";
		(Bmult[11] => Cmult[31]) = "";
		(Bmult[12] => Cmult[31]) = "";
		(Bmult[13] => Cmult[31]) = "";
		(Bmult[14] => Cmult[31]) = "";
		(Bmult[15] => Cmult[31]) = "";
		(Bmult[16] => Cmult[31]) = "";
		(Bmult[17] => Cmult[31]) = "";
		(Bmult[18] => Cmult[31]) = "";
		(Bmult[19] => Cmult[31]) = "";
		(Bmult[20] => Cmult[31]) = "";
		(Bmult[21] => Cmult[31]) = "";
		(Bmult[22] => Cmult[31]) = "";
		(Bmult[23] => Cmult[31]) = "";
		(Bmult[24] => Cmult[31]) = "";
		(Bmult[25] => Cmult[31]) = "";
		(Bmult[26] => Cmult[31]) = "";
		(Bmult[27] => Cmult[31]) = "";
		(Bmult[28] => Cmult[31]) = "";
		(Bmult[29] => Cmult[31]) = "";
		(Bmult[30] => Cmult[31]) = "";
		(Bmult[31] => Cmult[31]) = "";		
		(Valid_mult[0] => Cmult[31]) = "";
		(Valid_mult[1] => Cmult[31]) = "";
		(sel_mul_32x32 => Cmult[31]) = "";
		(Amult[0]  => Cmult[32]) = "";
		(Amult[1]  => Cmult[32]) = "";
		(Amult[2]  => Cmult[32]) = "";
		(Amult[3]  => Cmult[32]) = "";
		(Amult[4]  => Cmult[32]) = "";
		(Amult[5]  => Cmult[32]) = "";
		(Amult[6]  => Cmult[32]) = "";
		(Amult[7]  => Cmult[32]) = "";
		(Amult[8]  => Cmult[32]) = "";
		(Amult[9]  => Cmult[32]) = "";
		(Amult[10] => Cmult[32]) = "";
		(Amult[11] => Cmult[32]) = "";
		(Amult[12] => Cmult[32]) = "";
		(Amult[13] => Cmult[32]) = "";
		(Amult[14] => Cmult[32]) = "";
		(Amult[15] => Cmult[32]) = "";
		(Amult[16] => Cmult[32]) = "";
		(Amult[17] => Cmult[32]) = "";
		(Amult[18] => Cmult[32]) = "";
		(Amult[19] => Cmult[32]) = "";
		(Amult[20] => Cmult[32]) = "";
		(Amult[21] => Cmult[32]) = "";
		(Amult[22] => Cmult[32]) = "";
		(Amult[23] => Cmult[32]) = "";
		(Amult[24] => Cmult[32]) = "";
		(Amult[25] => Cmult[32]) = "";
		(Amult[26] => Cmult[32]) = "";
		(Amult[27] => Cmult[32]) = "";
		(Amult[28] => Cmult[32]) = "";
		(Amult[29] => Cmult[32]) = "";
		(Amult[30] => Cmult[32]) = "";
		(Amult[31] => Cmult[32]) = "";
		(Bmult[0]  => Cmult[32]) = "";
		(Bmult[1]  => Cmult[32]) = "";
		(Bmult[2]  => Cmult[32]) = "";
		(Bmult[3]  => Cmult[32]) = "";
		(Bmult[4]  => Cmult[32]) = "";
		(Bmult[5]  => Cmult[32]) = "";
		(Bmult[6]  => Cmult[32]) = "";
		(Bmult[7]  => Cmult[32]) = "";
		(Bmult[8]  => Cmult[32]) = "";
		(Bmult[9]  => Cmult[32]) = "";
		(Bmult[10] => Cmult[32]) = "";
		(Bmult[11] => Cmult[32]) = "";
		(Bmult[12] => Cmult[32]) = "";
		(Bmult[13] => Cmult[32]) = "";
		(Bmult[14] => Cmult[32]) = "";
		(Bmult[15] => Cmult[32]) = "";
		(Bmult[16] => Cmult[32]) = "";
		(Bmult[17] => Cmult[32]) = "";
		(Bmult[18] => Cmult[32]) = "";
		(Bmult[19] => Cmult[32]) = "";
		(Bmult[20] => Cmult[32]) = "";
		(Bmult[21] => Cmult[32]) = "";
		(Bmult[22] => Cmult[32]) = "";
		(Bmult[23] => Cmult[32]) = "";
		(Bmult[24] => Cmult[32]) = "";
		(Bmult[25] => Cmult[32]) = "";
		(Bmult[26] => Cmult[32]) = "";
		(Bmult[27] => Cmult[32]) = "";
		(Bmult[28] => Cmult[32]) = "";
		(Bmult[29] => Cmult[32]) = "";
		(Bmult[30] => Cmult[32]) = "";
		(Bmult[31] => Cmult[32]) = "";		
		(Valid_mult[0] => Cmult[32]) = "";
		(Valid_mult[1] => Cmult[32]) = "";
		(sel_mul_32x32 => Cmult[32]) = "";
		(Amult[0]  => Cmult[33]) = "";
		(Amult[1]  => Cmult[33]) = "";
		(Amult[2]  => Cmult[33]) = "";
		(Amult[3]  => Cmult[33]) = "";
		(Amult[4]  => Cmult[33]) = "";
		(Amult[5]  => Cmult[33]) = "";
		(Amult[6]  => Cmult[33]) = "";
		(Amult[7]  => Cmult[33]) = "";
		(Amult[8]  => Cmult[33]) = "";
		(Amult[9]  => Cmult[33]) = "";
		(Amult[10] => Cmult[33]) = "";
		(Amult[11] => Cmult[33]) = "";
		(Amult[12] => Cmult[33]) = "";
		(Amult[13] => Cmult[33]) = "";
		(Amult[14] => Cmult[33]) = "";
		(Amult[15] => Cmult[33]) = "";
		(Amult[16] => Cmult[33]) = "";
		(Amult[17] => Cmult[33]) = "";
		(Amult[18] => Cmult[33]) = "";
		(Amult[19] => Cmult[33]) = "";
		(Amult[20] => Cmult[33]) = "";
		(Amult[21] => Cmult[33]) = "";
		(Amult[22] => Cmult[33]) = "";
		(Amult[23] => Cmult[33]) = "";
		(Amult[24] => Cmult[33]) = "";
		(Amult[25] => Cmult[33]) = "";
		(Amult[26] => Cmult[33]) = "";
		(Amult[27] => Cmult[33]) = "";
		(Amult[28] => Cmult[33]) = "";
		(Amult[29] => Cmult[33]) = "";
		(Amult[30] => Cmult[33]) = "";
		(Amult[31] => Cmult[33]) = "";
		(Bmult[0]  => Cmult[33]) = "";
		(Bmult[1]  => Cmult[33]) = "";
		(Bmult[2]  => Cmult[33]) = "";
		(Bmult[3]  => Cmult[33]) = "";
		(Bmult[4]  => Cmult[33]) = "";
		(Bmult[5]  => Cmult[33]) = "";
		(Bmult[6]  => Cmult[33]) = "";
		(Bmult[7]  => Cmult[33]) = "";
		(Bmult[8]  => Cmult[33]) = "";
		(Bmult[9]  => Cmult[33]) = "";
		(Bmult[10] => Cmult[33]) = "";
		(Bmult[11] => Cmult[33]) = "";
		(Bmult[12] => Cmult[33]) = "";
		(Bmult[13] => Cmult[33]) = "";
		(Bmult[14] => Cmult[33]) = "";
		(Bmult[15] => Cmult[33]) = "";
		(Bmult[16] => Cmult[33]) = "";
		(Bmult[17] => Cmult[33]) = "";
		(Bmult[18] => Cmult[33]) = "";
		(Bmult[19] => Cmult[33]) = "";
		(Bmult[20] => Cmult[33]) = "";
		(Bmult[21] => Cmult[33]) = "";
		(Bmult[22] => Cmult[33]) = "";
		(Bmult[23] => Cmult[33]) = "";
		(Bmult[24] => Cmult[33]) = "";
		(Bmult[25] => Cmult[33]) = "";
		(Bmult[26] => Cmult[33]) = "";
		(Bmult[27] => Cmult[33]) = "";
		(Bmult[28] => Cmult[33]) = "";
		(Bmult[29] => Cmult[33]) = "";
		(Bmult[30] => Cmult[33]) = "";
		(Bmult[31] => Cmult[33]) = "";		
		(Valid_mult[0] => Cmult[33]) = "";
		(Valid_mult[1] => Cmult[33]) = "";
		(sel_mul_32x32 => Cmult[33]) = "";
		(Amult[0]  => Cmult[34]) = "";
		(Amult[1]  => Cmult[34]) = "";
		(Amult[2]  => Cmult[34]) = "";
		(Amult[3]  => Cmult[34]) = "";
		(Amult[4]  => Cmult[34]) = "";
		(Amult[5]  => Cmult[34]) = "";
		(Amult[6]  => Cmult[34]) = "";
		(Amult[7]  => Cmult[34]) = "";
		(Amult[8]  => Cmult[34]) = "";
		(Amult[9]  => Cmult[34]) = "";
		(Amult[10] => Cmult[34]) = "";
		(Amult[11] => Cmult[34]) = "";
		(Amult[12] => Cmult[34]) = "";
		(Amult[13] => Cmult[34]) = "";
		(Amult[14] => Cmult[34]) = "";
		(Amult[15] => Cmult[34]) = "";
		(Amult[16] => Cmult[34]) = "";
		(Amult[17] => Cmult[34]) = "";
		(Amult[18] => Cmult[34]) = "";
		(Amult[19] => Cmult[34]) = "";
		(Amult[20] => Cmult[34]) = "";
		(Amult[21] => Cmult[34]) = "";
		(Amult[22] => Cmult[34]) = "";
		(Amult[23] => Cmult[34]) = "";
		(Amult[24] => Cmult[34]) = "";
		(Amult[25] => Cmult[34]) = "";
		(Amult[26] => Cmult[34]) = "";
		(Amult[27] => Cmult[34]) = "";
		(Amult[28] => Cmult[34]) = "";
		(Amult[29] => Cmult[34]) = "";
		(Amult[30] => Cmult[34]) = "";
		(Amult[31] => Cmult[34]) = "";
		(Bmult[0]  => Cmult[34]) = "";
		(Bmult[1]  => Cmult[34]) = "";
		(Bmult[2]  => Cmult[34]) = "";
		(Bmult[3]  => Cmult[34]) = "";
		(Bmult[4]  => Cmult[34]) = "";
		(Bmult[5]  => Cmult[34]) = "";
		(Bmult[6]  => Cmult[34]) = "";
		(Bmult[7]  => Cmult[34]) = "";
		(Bmult[8]  => Cmult[34]) = "";
		(Bmult[9]  => Cmult[34]) = "";
		(Bmult[10] => Cmult[34]) = "";
		(Bmult[11] => Cmult[34]) = "";
		(Bmult[12] => Cmult[34]) = "";
		(Bmult[13] => Cmult[34]) = "";
		(Bmult[14] => Cmult[34]) = "";
		(Bmult[15] => Cmult[34]) = "";
		(Bmult[16] => Cmult[34]) = "";
		(Bmult[17] => Cmult[34]) = "";
		(Bmult[18] => Cmult[34]) = "";
		(Bmult[19] => Cmult[34]) = "";
		(Bmult[20] => Cmult[34]) = "";
		(Bmult[21] => Cmult[34]) = "";
		(Bmult[22] => Cmult[34]) = "";
		(Bmult[23] => Cmult[34]) = "";
		(Bmult[24] => Cmult[34]) = "";
		(Bmult[25] => Cmult[34]) = "";
		(Bmult[26] => Cmult[34]) = "";
		(Bmult[27] => Cmult[34]) = "";
		(Bmult[28] => Cmult[34]) = "";
		(Bmult[29] => Cmult[34]) = "";
		(Bmult[30] => Cmult[34]) = "";
		(Bmult[31] => Cmult[34]) = "";		
		(Valid_mult[0] => Cmult[34]) = "";
		(Valid_mult[1] => Cmult[34]) = "";
		(sel_mul_32x32 => Cmult[34]) = "";
		(Amult[0]  => Cmult[35]) = "";
		(Amult[1]  => Cmult[35]) = "";
		(Amult[2]  => Cmult[35]) = "";
		(Amult[3]  => Cmult[35]) = "";
		(Amult[4]  => Cmult[35]) = "";
		(Amult[5]  => Cmult[35]) = "";
		(Amult[6]  => Cmult[35]) = "";
		(Amult[7]  => Cmult[35]) = "";
		(Amult[8]  => Cmult[35]) = "";
		(Amult[9]  => Cmult[35]) = "";
		(Amult[10] => Cmult[35]) = "";
		(Amult[11] => Cmult[35]) = "";
		(Amult[12] => Cmult[35]) = "";
		(Amult[13] => Cmult[35]) = "";
		(Amult[14] => Cmult[35]) = "";
		(Amult[15] => Cmult[35]) = "";
		(Amult[16] => Cmult[35]) = "";
		(Amult[17] => Cmult[35]) = "";
		(Amult[18] => Cmult[35]) = "";
		(Amult[19] => Cmult[35]) = "";
		(Amult[20] => Cmult[35]) = "";
		(Amult[21] => Cmult[35]) = "";
		(Amult[22] => Cmult[35]) = "";
		(Amult[23] => Cmult[35]) = "";
		(Amult[24] => Cmult[35]) = "";
		(Amult[25] => Cmult[35]) = "";
		(Amult[26] => Cmult[35]) = "";
		(Amult[27] => Cmult[35]) = "";
		(Amult[28] => Cmult[35]) = "";
		(Amult[29] => Cmult[35]) = "";
		(Amult[30] => Cmult[35]) = "";
		(Amult[31] => Cmult[35]) = "";
		(Bmult[0]  => Cmult[35]) = "";
		(Bmult[1]  => Cmult[35]) = "";
		(Bmult[2]  => Cmult[35]) = "";
		(Bmult[3]  => Cmult[35]) = "";
		(Bmult[4]  => Cmult[35]) = "";
		(Bmult[5]  => Cmult[35]) = "";
		(Bmult[6]  => Cmult[35]) = "";
		(Bmult[7]  => Cmult[35]) = "";
		(Bmult[8]  => Cmult[35]) = "";
		(Bmult[9]  => Cmult[35]) = "";
		(Bmult[10] => Cmult[35]) = "";
		(Bmult[11] => Cmult[35]) = "";
		(Bmult[12] => Cmult[35]) = "";
		(Bmult[13] => Cmult[35]) = "";
		(Bmult[14] => Cmult[35]) = "";
		(Bmult[15] => Cmult[35]) = "";
		(Bmult[16] => Cmult[35]) = "";
		(Bmult[17] => Cmult[35]) = "";
		(Bmult[18] => Cmult[35]) = "";
		(Bmult[19] => Cmult[35]) = "";
		(Bmult[20] => Cmult[35]) = "";
		(Bmult[21] => Cmult[35]) = "";
		(Bmult[22] => Cmult[35]) = "";
		(Bmult[23] => Cmult[35]) = "";
		(Bmult[24] => Cmult[35]) = "";
		(Bmult[25] => Cmult[35]) = "";
		(Bmult[26] => Cmult[35]) = "";
		(Bmult[27] => Cmult[35]) = "";
		(Bmult[28] => Cmult[35]) = "";
		(Bmult[29] => Cmult[35]) = "";
		(Bmult[30] => Cmult[35]) = "";
		(Bmult[31] => Cmult[35]) = "";		
		(Valid_mult[0] => Cmult[35]) = "";
		(Valid_mult[1] => Cmult[35]) = "";
		(sel_mul_32x32 => Cmult[35]) = "";
		(Amult[0]  => Cmult[36]) = "";
		(Amult[1]  => Cmult[36]) = "";
		(Amult[2]  => Cmult[36]) = "";
		(Amult[3]  => Cmult[36]) = "";
		(Amult[4]  => Cmult[36]) = "";
		(Amult[5]  => Cmult[36]) = "";
		(Amult[6]  => Cmult[36]) = "";
		(Amult[7]  => Cmult[36]) = "";
		(Amult[8]  => Cmult[36]) = "";
		(Amult[9]  => Cmult[36]) = "";
		(Amult[10] => Cmult[36]) = "";
		(Amult[11] => Cmult[36]) = "";
		(Amult[12] => Cmult[36]) = "";
		(Amult[13] => Cmult[36]) = "";
		(Amult[14] => Cmult[36]) = "";
		(Amult[15] => Cmult[36]) = "";
		(Amult[16] => Cmult[36]) = "";
		(Amult[17] => Cmult[36]) = "";
		(Amult[18] => Cmult[36]) = "";
		(Amult[19] => Cmult[36]) = "";
		(Amult[20] => Cmult[36]) = "";
		(Amult[21] => Cmult[36]) = "";
		(Amult[22] => Cmult[36]) = "";
		(Amult[23] => Cmult[36]) = "";
		(Amult[24] => Cmult[36]) = "";
		(Amult[25] => Cmult[36]) = "";
		(Amult[26] => Cmult[36]) = "";
		(Amult[27] => Cmult[36]) = "";
		(Amult[28] => Cmult[36]) = "";
		(Amult[29] => Cmult[36]) = "";
		(Amult[30] => Cmult[36]) = "";
		(Amult[31] => Cmult[36]) = "";
		(Bmult[0]  => Cmult[36]) = "";
		(Bmult[1]  => Cmult[36]) = "";
		(Bmult[2]  => Cmult[36]) = "";
		(Bmult[3]  => Cmult[36]) = "";
		(Bmult[4]  => Cmult[36]) = "";
		(Bmult[5]  => Cmult[36]) = "";
		(Bmult[6]  => Cmult[36]) = "";
		(Bmult[7]  => Cmult[36]) = "";
		(Bmult[8]  => Cmult[36]) = "";
		(Bmult[9]  => Cmult[36]) = "";
		(Bmult[10] => Cmult[36]) = "";
		(Bmult[11] => Cmult[36]) = "";
		(Bmult[12] => Cmult[36]) = "";
		(Bmult[13] => Cmult[36]) = "";
		(Bmult[14] => Cmult[36]) = "";
		(Bmult[15] => Cmult[36]) = "";
		(Bmult[16] => Cmult[36]) = "";
		(Bmult[17] => Cmult[36]) = "";
		(Bmult[18] => Cmult[36]) = "";
		(Bmult[19] => Cmult[36]) = "";
		(Bmult[20] => Cmult[36]) = "";
		(Bmult[21] => Cmult[36]) = "";
		(Bmult[22] => Cmult[36]) = "";
		(Bmult[23] => Cmult[36]) = "";
		(Bmult[24] => Cmult[36]) = "";
		(Bmult[25] => Cmult[36]) = "";
		(Bmult[26] => Cmult[36]) = "";
		(Bmult[27] => Cmult[36]) = "";
		(Bmult[28] => Cmult[36]) = "";
		(Bmult[29] => Cmult[36]) = "";
		(Bmult[30] => Cmult[36]) = "";
		(Bmult[31] => Cmult[36]) = "";		
		(Valid_mult[0] => Cmult[36]) = "";
		(Valid_mult[1] => Cmult[36]) = "";
		(sel_mul_32x32 => Cmult[36]) = "";
		(Amult[0]  => Cmult[37]) = "";
		(Amult[1]  => Cmult[37]) = "";
		(Amult[2]  => Cmult[37]) = "";
		(Amult[3]  => Cmult[37]) = "";
		(Amult[4]  => Cmult[37]) = "";
		(Amult[5]  => Cmult[37]) = "";
		(Amult[6]  => Cmult[37]) = "";
		(Amult[7]  => Cmult[37]) = "";
		(Amult[8]  => Cmult[37]) = "";
		(Amult[9]  => Cmult[37]) = "";
		(Amult[10] => Cmult[37]) = "";
		(Amult[11] => Cmult[37]) = "";
		(Amult[12] => Cmult[37]) = "";
		(Amult[13] => Cmult[37]) = "";
		(Amult[14] => Cmult[37]) = "";
		(Amult[15] => Cmult[37]) = "";
		(Amult[16] => Cmult[37]) = "";
		(Amult[17] => Cmult[37]) = "";
		(Amult[18] => Cmult[37]) = "";
		(Amult[19] => Cmult[37]) = "";
		(Amult[20] => Cmult[37]) = "";
		(Amult[21] => Cmult[37]) = "";
		(Amult[22] => Cmult[37]) = "";
		(Amult[23] => Cmult[37]) = "";
		(Amult[24] => Cmult[37]) = "";
		(Amult[25] => Cmult[37]) = "";
		(Amult[26] => Cmult[37]) = "";
		(Amult[27] => Cmult[37]) = "";
		(Amult[28] => Cmult[37]) = "";
		(Amult[29] => Cmult[37]) = "";
		(Amult[30] => Cmult[37]) = "";
		(Amult[31] => Cmult[37]) = "";
		(Bmult[0]  => Cmult[37]) = "";
		(Bmult[1]  => Cmult[37]) = "";
		(Bmult[2]  => Cmult[37]) = "";
		(Bmult[3]  => Cmult[37]) = "";
		(Bmult[4]  => Cmult[37]) = "";
		(Bmult[5]  => Cmult[37]) = "";
		(Bmult[6]  => Cmult[37]) = "";
		(Bmult[7]  => Cmult[37]) = "";
		(Bmult[8]  => Cmult[37]) = "";
		(Bmult[9]  => Cmult[37]) = "";
		(Bmult[10] => Cmult[37]) = "";
		(Bmult[11] => Cmult[37]) = "";
		(Bmult[12] => Cmult[37]) = "";
		(Bmult[13] => Cmult[37]) = "";
		(Bmult[14] => Cmult[37]) = "";
		(Bmult[15] => Cmult[37]) = "";
		(Bmult[16] => Cmult[37]) = "";
		(Bmult[17] => Cmult[37]) = "";
		(Bmult[18] => Cmult[37]) = "";
		(Bmult[19] => Cmult[37]) = "";
		(Bmult[20] => Cmult[37]) = "";
		(Bmult[21] => Cmult[37]) = "";
		(Bmult[22] => Cmult[37]) = "";
		(Bmult[23] => Cmult[37]) = "";
		(Bmult[24] => Cmult[37]) = "";
		(Bmult[25] => Cmult[37]) = "";
		(Bmult[26] => Cmult[37]) = "";
		(Bmult[27] => Cmult[37]) = "";
		(Bmult[28] => Cmult[37]) = "";
		(Bmult[29] => Cmult[37]) = "";
		(Bmult[30] => Cmult[37]) = "";
		(Bmult[31] => Cmult[37]) = "";		
		(Valid_mult[0] => Cmult[37]) = "";
		(Valid_mult[1] => Cmult[37]) = "";
		(sel_mul_32x32 => Cmult[37]) = "";
		(Amult[0]  => Cmult[38]) = "";
		(Amult[1]  => Cmult[38]) = "";
		(Amult[2]  => Cmult[38]) = "";
		(Amult[3]  => Cmult[38]) = "";
		(Amult[4]  => Cmult[38]) = "";
		(Amult[5]  => Cmult[38]) = "";
		(Amult[6]  => Cmult[38]) = "";
		(Amult[7]  => Cmult[38]) = "";
		(Amult[8]  => Cmult[38]) = "";
		(Amult[9]  => Cmult[38]) = "";
		(Amult[10] => Cmult[38]) = "";
		(Amult[11] => Cmult[38]) = "";
		(Amult[12] => Cmult[38]) = "";
		(Amult[13] => Cmult[38]) = "";
		(Amult[14] => Cmult[38]) = "";
		(Amult[15] => Cmult[38]) = "";
		(Amult[16] => Cmult[38]) = "";
		(Amult[17] => Cmult[38]) = "";
		(Amult[18] => Cmult[38]) = "";
		(Amult[19] => Cmult[38]) = "";
		(Amult[20] => Cmult[38]) = "";
		(Amult[21] => Cmult[38]) = "";
		(Amult[22] => Cmult[38]) = "";
		(Amult[23] => Cmult[38]) = "";
		(Amult[24] => Cmult[38]) = "";
		(Amult[25] => Cmult[38]) = "";
		(Amult[26] => Cmult[38]) = "";
		(Amult[27] => Cmult[38]) = "";
		(Amult[28] => Cmult[38]) = "";
		(Amult[29] => Cmult[38]) = "";
		(Amult[30] => Cmult[38]) = "";
		(Amult[31] => Cmult[38]) = "";
		(Bmult[0]  => Cmult[38]) = "";
		(Bmult[1]  => Cmult[38]) = "";
		(Bmult[2]  => Cmult[38]) = "";
		(Bmult[3]  => Cmult[38]) = "";
		(Bmult[4]  => Cmult[38]) = "";
		(Bmult[5]  => Cmult[38]) = "";
		(Bmult[6]  => Cmult[38]) = "";
		(Bmult[7]  => Cmult[38]) = "";
		(Bmult[8]  => Cmult[38]) = "";
		(Bmult[9]  => Cmult[38]) = "";
		(Bmult[10] => Cmult[38]) = "";
		(Bmult[11] => Cmult[38]) = "";
		(Bmult[12] => Cmult[38]) = "";
		(Bmult[13] => Cmult[38]) = "";
		(Bmult[14] => Cmult[38]) = "";
		(Bmult[15] => Cmult[38]) = "";
		(Bmult[16] => Cmult[38]) = "";
		(Bmult[17] => Cmult[38]) = "";
		(Bmult[18] => Cmult[38]) = "";
		(Bmult[19] => Cmult[38]) = "";
		(Bmult[20] => Cmult[38]) = "";
		(Bmult[21] => Cmult[38]) = "";
		(Bmult[22] => Cmult[38]) = "";
		(Bmult[23] => Cmult[38]) = "";
		(Bmult[24] => Cmult[38]) = "";
		(Bmult[25] => Cmult[38]) = "";
		(Bmult[26] => Cmult[38]) = "";
		(Bmult[27] => Cmult[38]) = "";
		(Bmult[28] => Cmult[38]) = "";
		(Bmult[29] => Cmult[38]) = "";
		(Bmult[30] => Cmult[38]) = "";
		(Bmult[31] => Cmult[38]) = "";		
		(Valid_mult[0] => Cmult[38]) = "";
		(Valid_mult[1] => Cmult[38]) = "";
		(sel_mul_32x32 => Cmult[38]) = "";	
		(Amult[0]  => Cmult[39]) = "";
		(Amult[1]  => Cmult[39]) = "";
		(Amult[2]  => Cmult[39]) = "";
		(Amult[3]  => Cmult[39]) = "";
		(Amult[4]  => Cmult[39]) = "";
		(Amult[5]  => Cmult[39]) = "";
		(Amult[6]  => Cmult[39]) = "";
		(Amult[7]  => Cmult[39]) = "";
		(Amult[8]  => Cmult[39]) = "";
		(Amult[9]  => Cmult[39]) = "";
		(Amult[10] => Cmult[39]) = "";
		(Amult[11] => Cmult[39]) = "";
		(Amult[12] => Cmult[39]) = "";
		(Amult[13] => Cmult[39]) = "";
		(Amult[14] => Cmult[39]) = "";
		(Amult[15] => Cmult[39]) = "";
		(Amult[16] => Cmult[39]) = "";
		(Amult[17] => Cmult[39]) = "";
		(Amult[18] => Cmult[39]) = "";
		(Amult[19] => Cmult[39]) = "";
		(Amult[20] => Cmult[39]) = "";
		(Amult[21] => Cmult[39]) = "";
		(Amult[22] => Cmult[39]) = "";
		(Amult[23] => Cmult[39]) = "";
		(Amult[24] => Cmult[39]) = "";
		(Amult[25] => Cmult[39]) = "";
		(Amult[26] => Cmult[39]) = "";
		(Amult[27] => Cmult[39]) = "";
		(Amult[28] => Cmult[39]) = "";
		(Amult[29] => Cmult[39]) = "";
		(Amult[30] => Cmult[39]) = "";
		(Amult[31] => Cmult[39]) = "";
		(Bmult[0]  => Cmult[39]) = "";
		(Bmult[1]  => Cmult[39]) = "";
		(Bmult[2]  => Cmult[39]) = "";
		(Bmult[3]  => Cmult[39]) = "";
		(Bmult[4]  => Cmult[39]) = "";
		(Bmult[5]  => Cmult[39]) = "";
		(Bmult[6]  => Cmult[39]) = "";
		(Bmult[7]  => Cmult[39]) = "";
		(Bmult[8]  => Cmult[39]) = "";
		(Bmult[9]  => Cmult[39]) = "";
		(Bmult[10] => Cmult[39]) = "";
		(Bmult[11] => Cmult[39]) = "";
		(Bmult[12] => Cmult[39]) = "";
		(Bmult[13] => Cmult[39]) = "";
		(Bmult[14] => Cmult[39]) = "";
		(Bmult[15] => Cmult[39]) = "";
		(Bmult[16] => Cmult[39]) = "";
		(Bmult[17] => Cmult[39]) = "";
		(Bmult[18] => Cmult[39]) = "";
		(Bmult[19] => Cmult[39]) = "";
		(Bmult[20] => Cmult[39]) = "";
		(Bmult[21] => Cmult[39]) = "";
		(Bmult[22] => Cmult[39]) = "";
		(Bmult[23] => Cmult[39]) = "";
		(Bmult[24] => Cmult[39]) = "";
		(Bmult[25] => Cmult[39]) = "";
		(Bmult[26] => Cmult[39]) = "";
		(Bmult[27] => Cmult[39]) = "";
		(Bmult[28] => Cmult[39]) = "";
		(Bmult[29] => Cmult[39]) = "";
		(Bmult[30] => Cmult[39]) = "";
		(Bmult[31] => Cmult[39]) = "";		
		(Valid_mult[0] => Cmult[39]) = "";
		(Valid_mult[1] => Cmult[39]) = "";
		(sel_mul_32x32 => Cmult[39]) = "";
		(Amult[0]  => Cmult[40]) = "";
		(Amult[1]  => Cmult[40]) = "";
		(Amult[2]  => Cmult[40]) = "";
		(Amult[3]  => Cmult[40]) = "";
		(Amult[4]  => Cmult[40]) = "";
		(Amult[5]  => Cmult[40]) = "";
		(Amult[6]  => Cmult[40]) = "";
		(Amult[7]  => Cmult[40]) = "";
		(Amult[8]  => Cmult[40]) = "";
		(Amult[9]  => Cmult[40]) = "";
		(Amult[10] => Cmult[40]) = "";
		(Amult[11] => Cmult[40]) = "";
		(Amult[12] => Cmult[40]) = "";
		(Amult[13] => Cmult[40]) = "";
		(Amult[14] => Cmult[40]) = "";
		(Amult[15] => Cmult[40]) = "";
		(Amult[16] => Cmult[40]) = "";
		(Amult[17] => Cmult[40]) = "";
		(Amult[18] => Cmult[40]) = "";
		(Amult[19] => Cmult[40]) = "";
		(Amult[20] => Cmult[40]) = "";
		(Amult[21] => Cmult[40]) = "";
		(Amult[22] => Cmult[40]) = "";
		(Amult[23] => Cmult[40]) = "";
		(Amult[24] => Cmult[40]) = "";
		(Amult[25] => Cmult[40]) = "";
		(Amult[26] => Cmult[40]) = "";
		(Amult[27] => Cmult[40]) = "";
		(Amult[28] => Cmult[40]) = "";
		(Amult[29] => Cmult[40]) = "";
		(Amult[30] => Cmult[40]) = "";
		(Amult[31] => Cmult[40]) = "";
		(Bmult[0]  => Cmult[40]) = "";
		(Bmult[1]  => Cmult[40]) = "";
		(Bmult[2]  => Cmult[40]) = "";
		(Bmult[3]  => Cmult[40]) = "";
		(Bmult[4]  => Cmult[40]) = "";
		(Bmult[5]  => Cmult[40]) = "";
		(Bmult[6]  => Cmult[40]) = "";
		(Bmult[7]  => Cmult[40]) = "";
		(Bmult[8]  => Cmult[40]) = "";
		(Bmult[9]  => Cmult[40]) = "";
		(Bmult[10] => Cmult[40]) = "";
		(Bmult[11] => Cmult[40]) = "";
		(Bmult[12] => Cmult[40]) = "";
		(Bmult[13] => Cmult[40]) = "";
		(Bmult[14] => Cmult[40]) = "";
		(Bmult[15] => Cmult[40]) = "";
		(Bmult[16] => Cmult[40]) = "";
		(Bmult[17] => Cmult[40]) = "";
		(Bmult[18] => Cmult[40]) = "";
		(Bmult[19] => Cmult[40]) = "";
		(Bmult[20] => Cmult[40]) = "";
		(Bmult[21] => Cmult[40]) = "";
		(Bmult[22] => Cmult[40]) = "";
		(Bmult[23] => Cmult[40]) = "";
		(Bmult[24] => Cmult[40]) = "";
		(Bmult[25] => Cmult[40]) = "";
		(Bmult[26] => Cmult[40]) = "";
		(Bmult[27] => Cmult[40]) = "";
		(Bmult[28] => Cmult[40]) = "";
		(Bmult[29] => Cmult[40]) = "";
		(Bmult[30] => Cmult[40]) = "";
		(Bmult[31] => Cmult[40]) = "";		
		(Valid_mult[0] => Cmult[40]) = "";
		(Valid_mult[1] => Cmult[40]) = "";
		(sel_mul_32x32 => Cmult[40]) = "";
		(Amult[0]  => Cmult[41]) = "";
		(Amult[1]  => Cmult[41]) = "";
		(Amult[2]  => Cmult[41]) = "";
		(Amult[3]  => Cmult[41]) = "";
		(Amult[4]  => Cmult[41]) = "";
		(Amult[5]  => Cmult[41]) = "";
		(Amult[6]  => Cmult[41]) = "";
		(Amult[7]  => Cmult[41]) = "";
		(Amult[8]  => Cmult[41]) = "";
		(Amult[9]  => Cmult[41]) = "";
		(Amult[10] => Cmult[41]) = "";
		(Amult[11] => Cmult[41]) = "";
		(Amult[12] => Cmult[41]) = "";
		(Amult[13] => Cmult[41]) = "";
		(Amult[14] => Cmult[41]) = "";
		(Amult[15] => Cmult[41]) = "";
		(Amult[16] => Cmult[41]) = "";
		(Amult[17] => Cmult[41]) = "";
		(Amult[18] => Cmult[41]) = "";
		(Amult[19] => Cmult[41]) = "";
		(Amult[20] => Cmult[41]) = "";
		(Amult[21] => Cmult[41]) = "";
		(Amult[22] => Cmult[41]) = "";
		(Amult[23] => Cmult[41]) = "";
		(Amult[24] => Cmult[41]) = "";
		(Amult[25] => Cmult[41]) = "";
		(Amult[26] => Cmult[41]) = "";
		(Amult[27] => Cmult[41]) = "";
		(Amult[28] => Cmult[41]) = "";
		(Amult[29] => Cmult[41]) = "";
		(Amult[30] => Cmult[41]) = "";
		(Amult[31] => Cmult[41]) = "";
		(Bmult[0]  => Cmult[41]) = "";
		(Bmult[1]  => Cmult[41]) = "";
		(Bmult[2]  => Cmult[41]) = "";
		(Bmult[3]  => Cmult[41]) = "";
		(Bmult[4]  => Cmult[41]) = "";
		(Bmult[5]  => Cmult[41]) = "";
		(Bmult[6]  => Cmult[41]) = "";
		(Bmult[7]  => Cmult[41]) = "";
		(Bmult[8]  => Cmult[41]) = "";
		(Bmult[9]  => Cmult[41]) = "";
		(Bmult[10] => Cmult[41]) = "";
		(Bmult[11] => Cmult[41]) = "";
		(Bmult[12] => Cmult[41]) = "";
		(Bmult[13] => Cmult[41]) = "";
		(Bmult[14] => Cmult[41]) = "";
		(Bmult[15] => Cmult[41]) = "";
		(Bmult[16] => Cmult[41]) = "";
		(Bmult[17] => Cmult[41]) = "";
		(Bmult[18] => Cmult[41]) = "";
		(Bmult[19] => Cmult[41]) = "";
		(Bmult[20] => Cmult[41]) = "";
		(Bmult[21] => Cmult[41]) = "";
		(Bmult[22] => Cmult[41]) = "";
		(Bmult[23] => Cmult[41]) = "";
		(Bmult[24] => Cmult[41]) = "";
		(Bmult[25] => Cmult[41]) = "";
		(Bmult[26] => Cmult[41]) = "";
		(Bmult[27] => Cmult[41]) = "";
		(Bmult[28] => Cmult[41]) = "";
		(Bmult[29] => Cmult[41]) = "";
		(Bmult[30] => Cmult[41]) = "";
		(Bmult[31] => Cmult[41]) = "";		
		(Valid_mult[0] => Cmult[41]) = "";
		(Valid_mult[1] => Cmult[41]) = "";
		(sel_mul_32x32 => Cmult[41]) = "";
		(Amult[0]  => Cmult[42]) = "";
		(Amult[1]  => Cmult[42]) = "";
		(Amult[2]  => Cmult[42]) = "";
		(Amult[3]  => Cmult[42]) = "";
		(Amult[4]  => Cmult[42]) = "";
		(Amult[5]  => Cmult[42]) = "";
		(Amult[6]  => Cmult[42]) = "";
		(Amult[7]  => Cmult[42]) = "";
		(Amult[8]  => Cmult[42]) = "";
		(Amult[9]  => Cmult[42]) = "";
		(Amult[10] => Cmult[42]) = "";
		(Amult[11] => Cmult[42]) = "";
		(Amult[12] => Cmult[42]) = "";
		(Amult[13] => Cmult[42]) = "";
		(Amult[14] => Cmult[42]) = "";
		(Amult[15] => Cmult[42]) = "";
		(Amult[16] => Cmult[42]) = "";
		(Amult[17] => Cmult[42]) = "";
		(Amult[18] => Cmult[42]) = "";
		(Amult[19] => Cmult[42]) = "";
		(Amult[20] => Cmult[42]) = "";
		(Amult[21] => Cmult[42]) = "";
		(Amult[22] => Cmult[42]) = "";
		(Amult[23] => Cmult[42]) = "";
		(Amult[24] => Cmult[42]) = "";
		(Amult[25] => Cmult[42]) = "";
		(Amult[26] => Cmult[42]) = "";
		(Amult[27] => Cmult[42]) = "";
		(Amult[28] => Cmult[42]) = "";
		(Amult[29] => Cmult[42]) = "";
		(Amult[30] => Cmult[42]) = "";
		(Amult[31] => Cmult[42]) = "";
		(Bmult[0]  => Cmult[42]) = "";
		(Bmult[1]  => Cmult[42]) = "";
		(Bmult[2]  => Cmult[42]) = "";
		(Bmult[3]  => Cmult[42]) = "";
		(Bmult[4]  => Cmult[42]) = "";
		(Bmult[5]  => Cmult[42]) = "";
		(Bmult[6]  => Cmult[42]) = "";
		(Bmult[7]  => Cmult[42]) = "";
		(Bmult[8]  => Cmult[42]) = "";
		(Bmult[9]  => Cmult[42]) = "";
		(Bmult[10] => Cmult[42]) = "";
		(Bmult[11] => Cmult[42]) = "";
		(Bmult[12] => Cmult[42]) = "";
		(Bmult[13] => Cmult[42]) = "";
		(Bmult[14] => Cmult[42]) = "";
		(Bmult[15] => Cmult[42]) = "";
		(Bmult[16] => Cmult[42]) = "";
		(Bmult[17] => Cmult[42]) = "";
		(Bmult[18] => Cmult[42]) = "";
		(Bmult[19] => Cmult[42]) = "";
		(Bmult[20] => Cmult[42]) = "";
		(Bmult[21] => Cmult[42]) = "";
		(Bmult[22] => Cmult[42]) = "";
		(Bmult[23] => Cmult[42]) = "";
		(Bmult[24] => Cmult[42]) = "";
		(Bmult[25] => Cmult[42]) = "";
		(Bmult[26] => Cmult[42]) = "";
		(Bmult[27] => Cmult[42]) = "";
		(Bmult[28] => Cmult[42]) = "";
		(Bmult[29] => Cmult[42]) = "";
		(Bmult[30] => Cmult[42]) = "";
		(Bmult[31] => Cmult[42]) = "";		
		(Valid_mult[0] => Cmult[42]) = "";
		(Valid_mult[1] => Cmult[42]) = "";
		(sel_mul_32x32 => Cmult[42]) = "";
		(Amult[0]  => Cmult[43]) = "";
		(Amult[1]  => Cmult[43]) = "";
		(Amult[2]  => Cmult[43]) = "";
		(Amult[3]  => Cmult[43]) = "";
		(Amult[4]  => Cmult[43]) = "";
		(Amult[5]  => Cmult[43]) = "";
		(Amult[6]  => Cmult[43]) = "";
		(Amult[7]  => Cmult[43]) = "";
		(Amult[8]  => Cmult[43]) = "";
		(Amult[9]  => Cmult[43]) = "";
		(Amult[10] => Cmult[43]) = "";
		(Amult[11] => Cmult[43]) = "";
		(Amult[12] => Cmult[43]) = "";
		(Amult[13] => Cmult[43]) = "";
		(Amult[14] => Cmult[43]) = "";
		(Amult[15] => Cmult[43]) = "";
		(Amult[16] => Cmult[43]) = "";
		(Amult[17] => Cmult[43]) = "";
		(Amult[18] => Cmult[43]) = "";
		(Amult[19] => Cmult[43]) = "";
		(Amult[20] => Cmult[43]) = "";
		(Amult[21] => Cmult[43]) = "";
		(Amult[22] => Cmult[43]) = "";
		(Amult[23] => Cmult[43]) = "";
		(Amult[24] => Cmult[43]) = "";
		(Amult[25] => Cmult[43]) = "";
		(Amult[26] => Cmult[43]) = "";
		(Amult[27] => Cmult[43]) = "";
		(Amult[28] => Cmult[43]) = "";
		(Amult[29] => Cmult[43]) = "";
		(Amult[30] => Cmult[43]) = "";
		(Amult[31] => Cmult[43]) = "";
		(Bmult[0]  => Cmult[43]) = "";
		(Bmult[1]  => Cmult[43]) = "";
		(Bmult[2]  => Cmult[43]) = "";
		(Bmult[3]  => Cmult[43]) = "";
		(Bmult[4]  => Cmult[43]) = "";
		(Bmult[5]  => Cmult[43]) = "";
		(Bmult[6]  => Cmult[43]) = "";
		(Bmult[7]  => Cmult[43]) = "";
		(Bmult[8]  => Cmult[43]) = "";
		(Bmult[9]  => Cmult[43]) = "";
		(Bmult[10] => Cmult[43]) = "";
		(Bmult[11] => Cmult[43]) = "";
		(Bmult[12] => Cmult[43]) = "";
		(Bmult[13] => Cmult[43]) = "";
		(Bmult[14] => Cmult[43]) = "";
		(Bmult[15] => Cmult[43]) = "";
		(Bmult[16] => Cmult[43]) = "";
		(Bmult[17] => Cmult[43]) = "";
		(Bmult[18] => Cmult[43]) = "";
		(Bmult[19] => Cmult[43]) = "";
		(Bmult[20] => Cmult[43]) = "";
		(Bmult[21] => Cmult[43]) = "";
		(Bmult[22] => Cmult[43]) = "";
		(Bmult[23] => Cmult[43]) = "";
		(Bmult[24] => Cmult[43]) = "";
		(Bmult[25] => Cmult[43]) = "";
		(Bmult[26] => Cmult[43]) = "";
		(Bmult[27] => Cmult[43]) = "";
		(Bmult[28] => Cmult[43]) = "";
		(Bmult[29] => Cmult[43]) = "";
		(Bmult[30] => Cmult[43]) = "";
		(Bmult[31] => Cmult[43]) = "";		
		(Valid_mult[0] => Cmult[43]) = "";
		(Valid_mult[1] => Cmult[43]) = "";
		(sel_mul_32x32 => Cmult[43]) = "";
		(Amult[0]  => Cmult[44]) = "";
		(Amult[1]  => Cmult[44]) = "";
		(Amult[2]  => Cmult[44]) = "";
		(Amult[3]  => Cmult[44]) = "";
		(Amult[4]  => Cmult[44]) = "";
		(Amult[5]  => Cmult[44]) = "";
		(Amult[6]  => Cmult[44]) = "";
		(Amult[7]  => Cmult[44]) = "";
		(Amult[8]  => Cmult[44]) = "";
		(Amult[9]  => Cmult[44]) = "";
		(Amult[10] => Cmult[44]) = "";
		(Amult[11] => Cmult[44]) = "";
		(Amult[12] => Cmult[44]) = "";
		(Amult[13] => Cmult[44]) = "";
		(Amult[14] => Cmult[44]) = "";
		(Amult[15] => Cmult[44]) = "";
		(Amult[16] => Cmult[44]) = "";
		(Amult[17] => Cmult[44]) = "";
		(Amult[18] => Cmult[44]) = "";
		(Amult[19] => Cmult[44]) = "";
		(Amult[20] => Cmult[44]) = "";
		(Amult[21] => Cmult[44]) = "";
		(Amult[22] => Cmult[44]) = "";
		(Amult[23] => Cmult[44]) = "";
		(Amult[24] => Cmult[44]) = "";
		(Amult[25] => Cmult[44]) = "";
		(Amult[26] => Cmult[44]) = "";
		(Amult[27] => Cmult[44]) = "";
		(Amult[28] => Cmult[44]) = "";
		(Amult[29] => Cmult[44]) = "";
		(Amult[30] => Cmult[44]) = "";
		(Amult[31] => Cmult[44]) = "";
		(Bmult[0]  => Cmult[44]) = "";
		(Bmult[1]  => Cmult[44]) = "";
		(Bmult[2]  => Cmult[44]) = "";
		(Bmult[3]  => Cmult[44]) = "";
		(Bmult[4]  => Cmult[44]) = "";
		(Bmult[5]  => Cmult[44]) = "";
		(Bmult[6]  => Cmult[44]) = "";
		(Bmult[7]  => Cmult[44]) = "";
		(Bmult[8]  => Cmult[44]) = "";
		(Bmult[9]  => Cmult[44]) = "";
		(Bmult[10] => Cmult[44]) = "";
		(Bmult[11] => Cmult[44]) = "";
		(Bmult[12] => Cmult[44]) = "";
		(Bmult[13] => Cmult[44]) = "";
		(Bmult[14] => Cmult[44]) = "";
		(Bmult[15] => Cmult[44]) = "";
		(Bmult[16] => Cmult[44]) = "";
		(Bmult[17] => Cmult[44]) = "";
		(Bmult[18] => Cmult[44]) = "";
		(Bmult[19] => Cmult[44]) = "";
		(Bmult[20] => Cmult[44]) = "";
		(Bmult[21] => Cmult[44]) = "";
		(Bmult[22] => Cmult[44]) = "";
		(Bmult[23] => Cmult[44]) = "";
		(Bmult[24] => Cmult[44]) = "";
		(Bmult[25] => Cmult[44]) = "";
		(Bmult[26] => Cmult[44]) = "";
		(Bmult[27] => Cmult[44]) = "";
		(Bmult[28] => Cmult[44]) = "";
		(Bmult[29] => Cmult[44]) = "";
		(Bmult[30] => Cmult[44]) = "";
		(Bmult[31] => Cmult[44]) = "";		
		(Valid_mult[0] => Cmult[44]) = "";
		(Valid_mult[1] => Cmult[44]) = "";
		(sel_mul_32x32 => Cmult[44]) = "";
		(Amult[0]  => Cmult[45]) = "";
		(Amult[1]  => Cmult[45]) = "";
		(Amult[2]  => Cmult[45]) = "";
		(Amult[3]  => Cmult[45]) = "";
		(Amult[4]  => Cmult[45]) = "";
		(Amult[5]  => Cmult[45]) = "";
		(Amult[6]  => Cmult[45]) = "";
		(Amult[7]  => Cmult[45]) = "";
		(Amult[8]  => Cmult[45]) = "";
		(Amult[9]  => Cmult[45]) = "";
		(Amult[10] => Cmult[45]) = "";
		(Amult[11] => Cmult[45]) = "";
		(Amult[12] => Cmult[45]) = "";
		(Amult[13] => Cmult[45]) = "";
		(Amult[14] => Cmult[45]) = "";
		(Amult[15] => Cmult[45]) = "";
		(Amult[16] => Cmult[45]) = "";
		(Amult[17] => Cmult[45]) = "";
		(Amult[18] => Cmult[45]) = "";
		(Amult[19] => Cmult[45]) = "";
		(Amult[20] => Cmult[45]) = "";
		(Amult[21] => Cmult[45]) = "";
		(Amult[22] => Cmult[45]) = "";
		(Amult[23] => Cmult[45]) = "";
		(Amult[24] => Cmult[45]) = "";
		(Amult[25] => Cmult[45]) = "";
		(Amult[26] => Cmult[45]) = "";
		(Amult[27] => Cmult[45]) = "";
		(Amult[28] => Cmult[45]) = "";
		(Amult[29] => Cmult[45]) = "";
		(Amult[30] => Cmult[45]) = "";
		(Amult[31] => Cmult[45]) = "";
		(Bmult[0]  => Cmult[45]) = "";
		(Bmult[1]  => Cmult[45]) = "";
		(Bmult[2]  => Cmult[45]) = "";
		(Bmult[3]  => Cmult[45]) = "";
		(Bmult[4]  => Cmult[45]) = "";
		(Bmult[5]  => Cmult[45]) = "";
		(Bmult[6]  => Cmult[45]) = "";
		(Bmult[7]  => Cmult[45]) = "";
		(Bmult[8]  => Cmult[45]) = "";
		(Bmult[9]  => Cmult[45]) = "";
		(Bmult[10] => Cmult[45]) = "";
		(Bmult[11] => Cmult[45]) = "";
		(Bmult[12] => Cmult[45]) = "";
		(Bmult[13] => Cmult[45]) = "";
		(Bmult[14] => Cmult[45]) = "";
		(Bmult[15] => Cmult[45]) = "";
		(Bmult[16] => Cmult[45]) = "";
		(Bmult[17] => Cmult[45]) = "";
		(Bmult[18] => Cmult[45]) = "";
		(Bmult[19] => Cmult[45]) = "";
		(Bmult[20] => Cmult[45]) = "";
		(Bmult[21] => Cmult[45]) = "";
		(Bmult[22] => Cmult[45]) = "";
		(Bmult[23] => Cmult[45]) = "";
		(Bmult[24] => Cmult[45]) = "";
		(Bmult[25] => Cmult[45]) = "";
		(Bmult[26] => Cmult[45]) = "";
		(Bmult[27] => Cmult[45]) = "";
		(Bmult[28] => Cmult[45]) = "";
		(Bmult[29] => Cmult[45]) = "";
		(Bmult[30] => Cmult[45]) = "";
		(Bmult[31] => Cmult[45]) = "";		
		(Valid_mult[0] => Cmult[45]) = "";
		(Valid_mult[1] => Cmult[45]) = "";
		(sel_mul_32x32 => Cmult[45]) = "";
		(Amult[0]  => Cmult[46]) = "";
		(Amult[1]  => Cmult[46]) = "";
		(Amult[2]  => Cmult[46]) = "";
		(Amult[3]  => Cmult[46]) = "";
		(Amult[4]  => Cmult[46]) = "";
		(Amult[5]  => Cmult[46]) = "";
		(Amult[6]  => Cmult[46]) = "";
		(Amult[7]  => Cmult[46]) = "";
		(Amult[8]  => Cmult[46]) = "";
		(Amult[9]  => Cmult[46]) = "";
		(Amult[10] => Cmult[46]) = "";
		(Amult[11] => Cmult[46]) = "";
		(Amult[12] => Cmult[46]) = "";
		(Amult[13] => Cmult[46]) = "";
		(Amult[14] => Cmult[46]) = "";
		(Amult[15] => Cmult[46]) = "";
		(Amult[16] => Cmult[46]) = "";
		(Amult[17] => Cmult[46]) = "";
		(Amult[18] => Cmult[46]) = "";
		(Amult[19] => Cmult[46]) = "";
		(Amult[20] => Cmult[46]) = "";
		(Amult[21] => Cmult[46]) = "";
		(Amult[22] => Cmult[46]) = "";
		(Amult[23] => Cmult[46]) = "";
		(Amult[24] => Cmult[46]) = "";
		(Amult[25] => Cmult[46]) = "";
		(Amult[26] => Cmult[46]) = "";
		(Amult[27] => Cmult[46]) = "";
		(Amult[28] => Cmult[46]) = "";
		(Amult[29] => Cmult[46]) = "";
		(Amult[30] => Cmult[46]) = "";
		(Amult[31] => Cmult[46]) = "";
		(Bmult[0]  => Cmult[46]) = "";
		(Bmult[1]  => Cmult[46]) = "";
		(Bmult[2]  => Cmult[46]) = "";
		(Bmult[3]  => Cmult[46]) = "";
		(Bmult[4]  => Cmult[46]) = "";
		(Bmult[5]  => Cmult[46]) = "";
		(Bmult[6]  => Cmult[46]) = "";
		(Bmult[7]  => Cmult[46]) = "";
		(Bmult[8]  => Cmult[46]) = "";
		(Bmult[9]  => Cmult[46]) = "";
		(Bmult[10] => Cmult[46]) = "";
		(Bmult[11] => Cmult[46]) = "";
		(Bmult[12] => Cmult[46]) = "";
		(Bmult[13] => Cmult[46]) = "";
		(Bmult[14] => Cmult[46]) = "";
		(Bmult[15] => Cmult[46]) = "";
		(Bmult[16] => Cmult[46]) = "";
		(Bmult[17] => Cmult[46]) = "";
		(Bmult[18] => Cmult[46]) = "";
		(Bmult[19] => Cmult[46]) = "";
		(Bmult[20] => Cmult[46]) = "";
		(Bmult[21] => Cmult[46]) = "";
		(Bmult[22] => Cmult[46]) = "";
		(Bmult[23] => Cmult[46]) = "";
		(Bmult[24] => Cmult[46]) = "";
		(Bmult[25] => Cmult[46]) = "";
		(Bmult[26] => Cmult[46]) = "";
		(Bmult[27] => Cmult[46]) = "";
		(Bmult[28] => Cmult[46]) = "";
		(Bmult[29] => Cmult[46]) = "";
		(Bmult[30] => Cmult[46]) = "";
		(Bmult[31] => Cmult[46]) = "";		
		(Valid_mult[0] => Cmult[46]) = "";
		(Valid_mult[1] => Cmult[46]) = "";
		(sel_mul_32x32 => Cmult[46]) = "";
		(Amult[0]  => Cmult[47]) = "";
		(Amult[1]  => Cmult[47]) = "";
		(Amult[2]  => Cmult[47]) = "";
		(Amult[3]  => Cmult[47]) = "";
		(Amult[4]  => Cmult[47]) = "";
		(Amult[5]  => Cmult[47]) = "";
		(Amult[6]  => Cmult[47]) = "";
		(Amult[7]  => Cmult[47]) = "";
		(Amult[8]  => Cmult[47]) = "";
		(Amult[9]  => Cmult[47]) = "";
		(Amult[10] => Cmult[47]) = "";
		(Amult[11] => Cmult[47]) = "";
		(Amult[12] => Cmult[47]) = "";
		(Amult[13] => Cmult[47]) = "";
		(Amult[14] => Cmult[47]) = "";
		(Amult[15] => Cmult[47]) = "";
		(Amult[16] => Cmult[47]) = "";
		(Amult[17] => Cmult[47]) = "";
		(Amult[18] => Cmult[47]) = "";
		(Amult[19] => Cmult[47]) = "";
		(Amult[20] => Cmult[47]) = "";
		(Amult[21] => Cmult[47]) = "";
		(Amult[22] => Cmult[47]) = "";
		(Amult[23] => Cmult[47]) = "";
		(Amult[24] => Cmult[47]) = "";
		(Amult[25] => Cmult[47]) = "";
		(Amult[26] => Cmult[47]) = "";
		(Amult[27] => Cmult[47]) = "";
		(Amult[28] => Cmult[47]) = "";
		(Amult[29] => Cmult[47]) = "";
		(Amult[30] => Cmult[47]) = "";
		(Amult[31] => Cmult[47]) = "";
		(Bmult[0]  => Cmult[47]) = "";
		(Bmult[1]  => Cmult[47]) = "";
		(Bmult[2]  => Cmult[47]) = "";
		(Bmult[3]  => Cmult[47]) = "";
		(Bmult[4]  => Cmult[47]) = "";
		(Bmult[5]  => Cmult[47]) = "";
		(Bmult[6]  => Cmult[47]) = "";
		(Bmult[7]  => Cmult[47]) = "";
		(Bmult[8]  => Cmult[47]) = "";
		(Bmult[9]  => Cmult[47]) = "";
		(Bmult[10] => Cmult[47]) = "";
		(Bmult[11] => Cmult[47]) = "";
		(Bmult[12] => Cmult[47]) = "";
		(Bmult[13] => Cmult[47]) = "";
		(Bmult[14] => Cmult[47]) = "";
		(Bmult[15] => Cmult[47]) = "";
		(Bmult[16] => Cmult[47]) = "";
		(Bmult[17] => Cmult[47]) = "";
		(Bmult[18] => Cmult[47]) = "";
		(Bmult[19] => Cmult[47]) = "";
		(Bmult[20] => Cmult[47]) = "";
		(Bmult[21] => Cmult[47]) = "";
		(Bmult[22] => Cmult[47]) = "";
		(Bmult[23] => Cmult[47]) = "";
		(Bmult[24] => Cmult[47]) = "";
		(Bmult[25] => Cmult[47]) = "";
		(Bmult[26] => Cmult[47]) = "";
		(Bmult[27] => Cmult[47]) = "";
		(Bmult[28] => Cmult[47]) = "";
		(Bmult[29] => Cmult[47]) = "";
		(Bmult[30] => Cmult[47]) = "";
		(Bmult[31] => Cmult[47]) = "";		
		(Valid_mult[0] => Cmult[47]) = "";
		(Valid_mult[1] => Cmult[47]) = "";
		(sel_mul_32x32 => Cmult[47]) = "";
		(Amult[0]  => Cmult[48]) = "";
		(Amult[1]  => Cmult[48]) = "";
		(Amult[2]  => Cmult[48]) = "";
		(Amult[3]  => Cmult[48]) = "";
		(Amult[4]  => Cmult[48]) = "";
		(Amult[5]  => Cmult[48]) = "";
		(Amult[6]  => Cmult[48]) = "";
		(Amult[7]  => Cmult[48]) = "";
		(Amult[8]  => Cmult[48]) = "";
		(Amult[9]  => Cmult[48]) = "";
		(Amult[10] => Cmult[48]) = "";
		(Amult[11] => Cmult[48]) = "";
		(Amult[12] => Cmult[48]) = "";
		(Amult[13] => Cmult[48]) = "";
		(Amult[14] => Cmult[48]) = "";
		(Amult[15] => Cmult[48]) = "";
		(Amult[16] => Cmult[48]) = "";
		(Amult[17] => Cmult[48]) = "";
		(Amult[18] => Cmult[48]) = "";
		(Amult[19] => Cmult[48]) = "";
		(Amult[20] => Cmult[48]) = "";
		(Amult[21] => Cmult[48]) = "";
		(Amult[22] => Cmult[48]) = "";
		(Amult[23] => Cmult[48]) = "";
		(Amult[24] => Cmult[48]) = "";
		(Amult[25] => Cmult[48]) = "";
		(Amult[26] => Cmult[48]) = "";
		(Amult[27] => Cmult[48]) = "";
		(Amult[28] => Cmult[48]) = "";
		(Amult[29] => Cmult[48]) = "";
		(Amult[30] => Cmult[48]) = "";
		(Amult[31] => Cmult[48]) = "";
		(Bmult[0]  => Cmult[48]) = "";
		(Bmult[1]  => Cmult[48]) = "";
		(Bmult[2]  => Cmult[48]) = "";
		(Bmult[3]  => Cmult[48]) = "";
		(Bmult[4]  => Cmult[48]) = "";
		(Bmult[5]  => Cmult[48]) = "";
		(Bmult[6]  => Cmult[48]) = "";
		(Bmult[7]  => Cmult[48]) = "";
		(Bmult[8]  => Cmult[48]) = "";
		(Bmult[9]  => Cmult[48]) = "";
		(Bmult[10] => Cmult[48]) = "";
		(Bmult[11] => Cmult[48]) = "";
		(Bmult[12] => Cmult[48]) = "";
		(Bmult[13] => Cmult[48]) = "";
		(Bmult[14] => Cmult[48]) = "";
		(Bmult[15] => Cmult[48]) = "";
		(Bmult[16] => Cmult[48]) = "";
		(Bmult[17] => Cmult[48]) = "";
		(Bmult[18] => Cmult[48]) = "";
		(Bmult[19] => Cmult[48]) = "";
		(Bmult[20] => Cmult[48]) = "";
		(Bmult[21] => Cmult[48]) = "";
		(Bmult[22] => Cmult[48]) = "";
		(Bmult[23] => Cmult[48]) = "";
		(Bmult[24] => Cmult[48]) = "";
		(Bmult[25] => Cmult[48]) = "";
		(Bmult[26] => Cmult[48]) = "";
		(Bmult[27] => Cmult[48]) = "";
		(Bmult[28] => Cmult[48]) = "";
		(Bmult[29] => Cmult[48]) = "";
		(Bmult[30] => Cmult[48]) = "";
		(Bmult[31] => Cmult[48]) = "";		
		(Valid_mult[0] => Cmult[48]) = "";
		(Valid_mult[1] => Cmult[48]) = "";
		(sel_mul_32x32 => Cmult[48]) = "";	
		(Amult[0]  => Cmult[49]) = "";
		(Amult[1]  => Cmult[49]) = "";
		(Amult[2]  => Cmult[49]) = "";
		(Amult[3]  => Cmult[49]) = "";
		(Amult[4]  => Cmult[49]) = "";
		(Amult[5]  => Cmult[49]) = "";
		(Amult[6]  => Cmult[49]) = "";
		(Amult[7]  => Cmult[49]) = "";
		(Amult[8]  => Cmult[49]) = "";
		(Amult[9]  => Cmult[49]) = "";
		(Amult[10] => Cmult[49]) = "";
		(Amult[11] => Cmult[49]) = "";
		(Amult[12] => Cmult[49]) = "";
		(Amult[13] => Cmult[49]) = "";
		(Amult[14] => Cmult[49]) = "";
		(Amult[15] => Cmult[49]) = "";
		(Amult[16] => Cmult[49]) = "";
		(Amult[17] => Cmult[49]) = "";
		(Amult[18] => Cmult[49]) = "";
		(Amult[19] => Cmult[49]) = "";
		(Amult[20] => Cmult[49]) = "";
		(Amult[21] => Cmult[49]) = "";
		(Amult[22] => Cmult[49]) = "";
		(Amult[23] => Cmult[49]) = "";
		(Amult[24] => Cmult[49]) = "";
		(Amult[25] => Cmult[49]) = "";
		(Amult[26] => Cmult[49]) = "";
		(Amult[27] => Cmult[49]) = "";
		(Amult[28] => Cmult[49]) = "";
		(Amult[29] => Cmult[49]) = "";
		(Amult[30] => Cmult[49]) = "";
		(Amult[31] => Cmult[49]) = "";
		(Bmult[0]  => Cmult[49]) = "";
		(Bmult[1]  => Cmult[49]) = "";
		(Bmult[2]  => Cmult[49]) = "";
		(Bmult[3]  => Cmult[49]) = "";
		(Bmult[4]  => Cmult[49]) = "";
		(Bmult[5]  => Cmult[49]) = "";
		(Bmult[6]  => Cmult[49]) = "";
		(Bmult[7]  => Cmult[49]) = "";
		(Bmult[8]  => Cmult[49]) = "";
		(Bmult[9]  => Cmult[49]) = "";
		(Bmult[10] => Cmult[49]) = "";
		(Bmult[11] => Cmult[49]) = "";
		(Bmult[12] => Cmult[49]) = "";
		(Bmult[13] => Cmult[49]) = "";
		(Bmult[14] => Cmult[49]) = "";
		(Bmult[15] => Cmult[49]) = "";
		(Bmult[16] => Cmult[49]) = "";
		(Bmult[17] => Cmult[49]) = "";
		(Bmult[18] => Cmult[49]) = "";
		(Bmult[19] => Cmult[49]) = "";
		(Bmult[20] => Cmult[49]) = "";
		(Bmult[21] => Cmult[49]) = "";
		(Bmult[22] => Cmult[49]) = "";
		(Bmult[23] => Cmult[49]) = "";
		(Bmult[24] => Cmult[49]) = "";
		(Bmult[25] => Cmult[49]) = "";
		(Bmult[26] => Cmult[49]) = "";
		(Bmult[27] => Cmult[49]) = "";
		(Bmult[28] => Cmult[49]) = "";
		(Bmult[29] => Cmult[49]) = "";
		(Bmult[30] => Cmult[49]) = "";
		(Bmult[31] => Cmult[49]) = "";		
		(Valid_mult[0] => Cmult[49]) = "";
		(Valid_mult[1] => Cmult[49]) = "";
		(sel_mul_32x32 => Cmult[49]) = "";
		(Amult[0]  => Cmult[50]) = "";
		(Amult[1]  => Cmult[50]) = "";
		(Amult[2]  => Cmult[50]) = "";
		(Amult[3]  => Cmult[50]) = "";
		(Amult[4]  => Cmult[50]) = "";
		(Amult[5]  => Cmult[50]) = "";
		(Amult[6]  => Cmult[50]) = "";
		(Amult[7]  => Cmult[50]) = "";
		(Amult[8]  => Cmult[50]) = "";
		(Amult[9]  => Cmult[50]) = "";
		(Amult[10] => Cmult[50]) = "";
		(Amult[11] => Cmult[50]) = "";
		(Amult[12] => Cmult[50]) = "";
		(Amult[13] => Cmult[50]) = "";
		(Amult[14] => Cmult[50]) = "";
		(Amult[15] => Cmult[50]) = "";
		(Amult[16] => Cmult[50]) = "";
		(Amult[17] => Cmult[50]) = "";
		(Amult[18] => Cmult[50]) = "";
		(Amult[19] => Cmult[50]) = "";
		(Amult[20] => Cmult[50]) = "";
		(Amult[21] => Cmult[50]) = "";
		(Amult[22] => Cmult[50]) = "";
		(Amult[23] => Cmult[50]) = "";
		(Amult[24] => Cmult[50]) = "";
		(Amult[25] => Cmult[50]) = "";
		(Amult[26] => Cmult[50]) = "";
		(Amult[27] => Cmult[50]) = "";
		(Amult[28] => Cmult[50]) = "";
		(Amult[29] => Cmult[50]) = "";
		(Amult[30] => Cmult[50]) = "";
		(Amult[31] => Cmult[50]) = "";
		(Bmult[0]  => Cmult[50]) = "";
		(Bmult[1]  => Cmult[50]) = "";
		(Bmult[2]  => Cmult[50]) = "";
		(Bmult[3]  => Cmult[50]) = "";
		(Bmult[4]  => Cmult[50]) = "";
		(Bmult[5]  => Cmult[50]) = "";
		(Bmult[6]  => Cmult[50]) = "";
		(Bmult[7]  => Cmult[50]) = "";
		(Bmult[8]  => Cmult[50]) = "";
		(Bmult[9]  => Cmult[50]) = "";
		(Bmult[10] => Cmult[50]) = "";
		(Bmult[11] => Cmult[50]) = "";
		(Bmult[12] => Cmult[50]) = "";
		(Bmult[13] => Cmult[50]) = "";
		(Bmult[14] => Cmult[50]) = "";
		(Bmult[15] => Cmult[50]) = "";
		(Bmult[16] => Cmult[50]) = "";
		(Bmult[17] => Cmult[50]) = "";
		(Bmult[18] => Cmult[50]) = "";
		(Bmult[19] => Cmult[50]) = "";
		(Bmult[20] => Cmult[50]) = "";
		(Bmult[21] => Cmult[50]) = "";
		(Bmult[22] => Cmult[50]) = "";
		(Bmult[23] => Cmult[50]) = "";
		(Bmult[24] => Cmult[50]) = "";
		(Bmult[25] => Cmult[50]) = "";
		(Bmult[26] => Cmult[50]) = "";
		(Bmult[27] => Cmult[50]) = "";
		(Bmult[28] => Cmult[50]) = "";
		(Bmult[29] => Cmult[50]) = "";
		(Bmult[30] => Cmult[50]) = "";
		(Bmult[31] => Cmult[50]) = "";		
		(Valid_mult[0] => Cmult[50]) = "";
		(Valid_mult[1] => Cmult[50]) = "";
		(sel_mul_32x32 => Cmult[50]) = "";
		(Amult[0]  => Cmult[51]) = "";
		(Amult[1]  => Cmult[51]) = "";
		(Amult[2]  => Cmult[51]) = "";
		(Amult[3]  => Cmult[51]) = "";
		(Amult[4]  => Cmult[51]) = "";
		(Amult[5]  => Cmult[51]) = "";
		(Amult[6]  => Cmult[51]) = "";
		(Amult[7]  => Cmult[51]) = "";
		(Amult[8]  => Cmult[51]) = "";
		(Amult[9]  => Cmult[51]) = "";
		(Amult[10] => Cmult[51]) = "";
		(Amult[11] => Cmult[51]) = "";
		(Amult[12] => Cmult[51]) = "";
		(Amult[13] => Cmult[51]) = "";
		(Amult[14] => Cmult[51]) = "";
		(Amult[15] => Cmult[51]) = "";
		(Amult[16] => Cmult[51]) = "";
		(Amult[17] => Cmult[51]) = "";
		(Amult[18] => Cmult[51]) = "";
		(Amult[19] => Cmult[51]) = "";
		(Amult[20] => Cmult[51]) = "";
		(Amult[21] => Cmult[51]) = "";
		(Amult[22] => Cmult[51]) = "";
		(Amult[23] => Cmult[51]) = "";
		(Amult[24] => Cmult[51]) = "";
		(Amult[25] => Cmult[51]) = "";
		(Amult[26] => Cmult[51]) = "";
		(Amult[27] => Cmult[51]) = "";
		(Amult[28] => Cmult[51]) = "";
		(Amult[29] => Cmult[51]) = "";
		(Amult[30] => Cmult[51]) = "";
		(Amult[31] => Cmult[51]) = "";
		(Bmult[0]  => Cmult[51]) = "";
		(Bmult[1]  => Cmult[51]) = "";
		(Bmult[2]  => Cmult[51]) = "";
		(Bmult[3]  => Cmult[51]) = "";
		(Bmult[4]  => Cmult[51]) = "";
		(Bmult[5]  => Cmult[51]) = "";
		(Bmult[6]  => Cmult[51]) = "";
		(Bmult[7]  => Cmult[51]) = "";
		(Bmult[8]  => Cmult[51]) = "";
		(Bmult[9]  => Cmult[51]) = "";
		(Bmult[10] => Cmult[51]) = "";
		(Bmult[11] => Cmult[51]) = "";
		(Bmult[12] => Cmult[51]) = "";
		(Bmult[13] => Cmult[51]) = "";
		(Bmult[14] => Cmult[51]) = "";
		(Bmult[15] => Cmult[51]) = "";
		(Bmult[16] => Cmult[51]) = "";
		(Bmult[17] => Cmult[51]) = "";
		(Bmult[18] => Cmult[51]) = "";
		(Bmult[19] => Cmult[51]) = "";
		(Bmult[20] => Cmult[51]) = "";
		(Bmult[21] => Cmult[51]) = "";
		(Bmult[22] => Cmult[51]) = "";
		(Bmult[23] => Cmult[51]) = "";
		(Bmult[24] => Cmult[51]) = "";
		(Bmult[25] => Cmult[51]) = "";
		(Bmult[26] => Cmult[51]) = "";
		(Bmult[27] => Cmult[51]) = "";
		(Bmult[28] => Cmult[51]) = "";
		(Bmult[29] => Cmult[51]) = "";
		(Bmult[30] => Cmult[51]) = "";
		(Bmult[31] => Cmult[51]) = "";		
		(Valid_mult[0] => Cmult[51]) = "";
		(Valid_mult[1] => Cmult[51]) = "";
		(sel_mul_32x32 => Cmult[51]) = "";
		(Amult[0]  => Cmult[52]) = "";
		(Amult[1]  => Cmult[52]) = "";
		(Amult[2]  => Cmult[52]) = "";
		(Amult[3]  => Cmult[52]) = "";
		(Amult[4]  => Cmult[52]) = "";
		(Amult[5]  => Cmult[52]) = "";
		(Amult[6]  => Cmult[52]) = "";
		(Amult[7]  => Cmult[52]) = "";
		(Amult[8]  => Cmult[52]) = "";
		(Amult[9]  => Cmult[52]) = "";
		(Amult[10] => Cmult[52]) = "";
		(Amult[11] => Cmult[52]) = "";
		(Amult[12] => Cmult[52]) = "";
		(Amult[13] => Cmult[52]) = "";
		(Amult[14] => Cmult[52]) = "";
		(Amult[15] => Cmult[52]) = "";
		(Amult[16] => Cmult[52]) = "";
		(Amult[17] => Cmult[52]) = "";
		(Amult[18] => Cmult[52]) = "";
		(Amult[19] => Cmult[52]) = "";
		(Amult[20] => Cmult[52]) = "";
		(Amult[21] => Cmult[52]) = "";
		(Amult[22] => Cmult[52]) = "";
		(Amult[23] => Cmult[52]) = "";
		(Amult[24] => Cmult[52]) = "";
		(Amult[25] => Cmult[52]) = "";
		(Amult[26] => Cmult[52]) = "";
		(Amult[27] => Cmult[52]) = "";
		(Amult[28] => Cmult[52]) = "";
		(Amult[29] => Cmult[52]) = "";
		(Amult[30] => Cmult[52]) = "";
		(Amult[31] => Cmult[52]) = "";
		(Bmult[0]  => Cmult[52]) = "";
		(Bmult[1]  => Cmult[52]) = "";
		(Bmult[2]  => Cmult[52]) = "";
		(Bmult[3]  => Cmult[52]) = "";
		(Bmult[4]  => Cmult[52]) = "";
		(Bmult[5]  => Cmult[52]) = "";
		(Bmult[6]  => Cmult[52]) = "";
		(Bmult[7]  => Cmult[52]) = "";
		(Bmult[8]  => Cmult[52]) = "";
		(Bmult[9]  => Cmult[52]) = "";
		(Bmult[10] => Cmult[52]) = "";
		(Bmult[11] => Cmult[52]) = "";
		(Bmult[12] => Cmult[52]) = "";
		(Bmult[13] => Cmult[52]) = "";
		(Bmult[14] => Cmult[52]) = "";
		(Bmult[15] => Cmult[52]) = "";
		(Bmult[16] => Cmult[52]) = "";
		(Bmult[17] => Cmult[52]) = "";
		(Bmult[18] => Cmult[52]) = "";
		(Bmult[19] => Cmult[52]) = "";
		(Bmult[20] => Cmult[52]) = "";
		(Bmult[21] => Cmult[52]) = "";
		(Bmult[22] => Cmult[52]) = "";
		(Bmult[23] => Cmult[52]) = "";
		(Bmult[24] => Cmult[52]) = "";
		(Bmult[25] => Cmult[52]) = "";
		(Bmult[26] => Cmult[52]) = "";
		(Bmult[27] => Cmult[52]) = "";
		(Bmult[28] => Cmult[52]) = "";
		(Bmult[29] => Cmult[52]) = "";
		(Bmult[30] => Cmult[52]) = "";
		(Bmult[31] => Cmult[52]) = "";		
		(Valid_mult[0] => Cmult[52]) = "";
		(Valid_mult[1] => Cmult[52]) = "";
		(sel_mul_32x32 => Cmult[52]) = "";
		(Amult[0]  => Cmult[53]) = "";
		(Amult[1]  => Cmult[53]) = "";
		(Amult[2]  => Cmult[53]) = "";
		(Amult[3]  => Cmult[53]) = "";
		(Amult[4]  => Cmult[53]) = "";
		(Amult[5]  => Cmult[53]) = "";
		(Amult[6]  => Cmult[53]) = "";
		(Amult[7]  => Cmult[53]) = "";
		(Amult[8]  => Cmult[53]) = "";
		(Amult[9]  => Cmult[53]) = "";
		(Amult[10] => Cmult[53]) = "";
		(Amult[11] => Cmult[53]) = "";
		(Amult[12] => Cmult[53]) = "";
		(Amult[13] => Cmult[53]) = "";
		(Amult[14] => Cmult[53]) = "";
		(Amult[15] => Cmult[53]) = "";
		(Amult[16] => Cmult[53]) = "";
		(Amult[17] => Cmult[53]) = "";
		(Amult[18] => Cmult[53]) = "";
		(Amult[19] => Cmult[53]) = "";
		(Amult[20] => Cmult[53]) = "";
		(Amult[21] => Cmult[53]) = "";
		(Amult[22] => Cmult[53]) = "";
		(Amult[23] => Cmult[53]) = "";
		(Amult[24] => Cmult[53]) = "";
		(Amult[25] => Cmult[53]) = "";
		(Amult[26] => Cmult[53]) = "";
		(Amult[27] => Cmult[53]) = "";
		(Amult[28] => Cmult[53]) = "";
		(Amult[29] => Cmult[53]) = "";
		(Amult[30] => Cmult[53]) = "";
		(Amult[31] => Cmult[53]) = "";
		(Bmult[0]  => Cmult[53]) = "";
		(Bmult[1]  => Cmult[53]) = "";
		(Bmult[2]  => Cmult[53]) = "";
		(Bmult[3]  => Cmult[53]) = "";
		(Bmult[4]  => Cmult[53]) = "";
		(Bmult[5]  => Cmult[53]) = "";
		(Bmult[6]  => Cmult[53]) = "";
		(Bmult[7]  => Cmult[53]) = "";
		(Bmult[8]  => Cmult[53]) = "";
		(Bmult[9]  => Cmult[53]) = "";
		(Bmult[10] => Cmult[53]) = "";
		(Bmult[11] => Cmult[53]) = "";
		(Bmult[12] => Cmult[53]) = "";
		(Bmult[13] => Cmult[53]) = "";
		(Bmult[14] => Cmult[53]) = "";
		(Bmult[15] => Cmult[53]) = "";
		(Bmult[16] => Cmult[53]) = "";
		(Bmult[17] => Cmult[53]) = "";
		(Bmult[18] => Cmult[53]) = "";
		(Bmult[19] => Cmult[53]) = "";
		(Bmult[20] => Cmult[53]) = "";
		(Bmult[21] => Cmult[53]) = "";
		(Bmult[22] => Cmult[53]) = "";
		(Bmult[23] => Cmult[53]) = "";
		(Bmult[24] => Cmult[53]) = "";
		(Bmult[25] => Cmult[53]) = "";
		(Bmult[26] => Cmult[53]) = "";
		(Bmult[27] => Cmult[53]) = "";
		(Bmult[28] => Cmult[53]) = "";
		(Bmult[29] => Cmult[53]) = "";
		(Bmult[30] => Cmult[53]) = "";
		(Bmult[31] => Cmult[53]) = "";		
		(Valid_mult[0] => Cmult[53]) = "";
		(Valid_mult[1] => Cmult[53]) = "";
		(sel_mul_32x32 => Cmult[53]) = "";
		(Amult[0]  => Cmult[54]) = "";
		(Amult[1]  => Cmult[54]) = "";
		(Amult[2]  => Cmult[54]) = "";
		(Amult[3]  => Cmult[54]) = "";
		(Amult[4]  => Cmult[54]) = "";
		(Amult[5]  => Cmult[54]) = "";
		(Amult[6]  => Cmult[54]) = "";
		(Amult[7]  => Cmult[54]) = "";
		(Amult[8]  => Cmult[54]) = "";
		(Amult[9]  => Cmult[54]) = "";
		(Amult[10] => Cmult[54]) = "";
		(Amult[11] => Cmult[54]) = "";
		(Amult[12] => Cmult[54]) = "";
		(Amult[13] => Cmult[54]) = "";
		(Amult[14] => Cmult[54]) = "";
		(Amult[15] => Cmult[54]) = "";
		(Amult[16] => Cmult[54]) = "";
		(Amult[17] => Cmult[54]) = "";
		(Amult[18] => Cmult[54]) = "";
		(Amult[19] => Cmult[54]) = "";
		(Amult[20] => Cmult[54]) = "";
		(Amult[21] => Cmult[54]) = "";
		(Amult[22] => Cmult[54]) = "";
		(Amult[23] => Cmult[54]) = "";
		(Amult[24] => Cmult[54]) = "";
		(Amult[25] => Cmult[54]) = "";
		(Amult[26] => Cmult[54]) = "";
		(Amult[27] => Cmult[54]) = "";
		(Amult[28] => Cmult[54]) = "";
		(Amult[29] => Cmult[54]) = "";
		(Amult[30] => Cmult[54]) = "";
		(Amult[31] => Cmult[54]) = "";
		(Bmult[0]  => Cmult[54]) = "";
		(Bmult[1]  => Cmult[54]) = "";
		(Bmult[2]  => Cmult[54]) = "";
		(Bmult[3]  => Cmult[54]) = "";
		(Bmult[4]  => Cmult[54]) = "";
		(Bmult[5]  => Cmult[54]) = "";
		(Bmult[6]  => Cmult[54]) = "";
		(Bmult[7]  => Cmult[54]) = "";
		(Bmult[8]  => Cmult[54]) = "";
		(Bmult[9]  => Cmult[54]) = "";
		(Bmult[10] => Cmult[54]) = "";
		(Bmult[11] => Cmult[54]) = "";
		(Bmult[12] => Cmult[54]) = "";
		(Bmult[13] => Cmult[54]) = "";
		(Bmult[14] => Cmult[54]) = "";
		(Bmult[15] => Cmult[54]) = "";
		(Bmult[16] => Cmult[54]) = "";
		(Bmult[17] => Cmult[54]) = "";
		(Bmult[18] => Cmult[54]) = "";
		(Bmult[19] => Cmult[54]) = "";
		(Bmult[20] => Cmult[54]) = "";
		(Bmult[21] => Cmult[54]) = "";
		(Bmult[22] => Cmult[54]) = "";
		(Bmult[23] => Cmult[54]) = "";
		(Bmult[24] => Cmult[54]) = "";
		(Bmult[25] => Cmult[54]) = "";
		(Bmult[26] => Cmult[54]) = "";
		(Bmult[27] => Cmult[54]) = "";
		(Bmult[28] => Cmult[54]) = "";
		(Bmult[29] => Cmult[54]) = "";
		(Bmult[30] => Cmult[54]) = "";
		(Bmult[31] => Cmult[54]) = "";		
		(Valid_mult[0] => Cmult[54]) = "";
		(Valid_mult[1] => Cmult[54]) = "";
		(sel_mul_32x32 => Cmult[54]) = "";
		(Amult[0]  => Cmult[55]) = "";
		(Amult[1]  => Cmult[55]) = "";
		(Amult[2]  => Cmult[55]) = "";
		(Amult[3]  => Cmult[55]) = "";
		(Amult[4]  => Cmult[55]) = "";
		(Amult[5]  => Cmult[55]) = "";
		(Amult[6]  => Cmult[55]) = "";
		(Amult[7]  => Cmult[55]) = "";
		(Amult[8]  => Cmult[55]) = "";
		(Amult[9]  => Cmult[55]) = "";
		(Amult[10] => Cmult[55]) = "";
		(Amult[11] => Cmult[55]) = "";
		(Amult[12] => Cmult[55]) = "";
		(Amult[13] => Cmult[55]) = "";
		(Amult[14] => Cmult[55]) = "";
		(Amult[15] => Cmult[55]) = "";
		(Amult[16] => Cmult[55]) = "";
		(Amult[17] => Cmult[55]) = "";
		(Amult[18] => Cmult[55]) = "";
		(Amult[19] => Cmult[55]) = "";
		(Amult[20] => Cmult[55]) = "";
		(Amult[21] => Cmult[55]) = "";
		(Amult[22] => Cmult[55]) = "";
		(Amult[23] => Cmult[55]) = "";
		(Amult[24] => Cmult[55]) = "";
		(Amult[25] => Cmult[55]) = "";
		(Amult[26] => Cmult[55]) = "";
		(Amult[27] => Cmult[55]) = "";
		(Amult[28] => Cmult[55]) = "";
		(Amult[29] => Cmult[55]) = "";
		(Amult[30] => Cmult[55]) = "";
		(Amult[31] => Cmult[55]) = "";
		(Bmult[0]  => Cmult[55]) = "";
		(Bmult[1]  => Cmult[55]) = "";
		(Bmult[2]  => Cmult[55]) = "";
		(Bmult[3]  => Cmult[55]) = "";
		(Bmult[4]  => Cmult[55]) = "";
		(Bmult[5]  => Cmult[55]) = "";
		(Bmult[6]  => Cmult[55]) = "";
		(Bmult[7]  => Cmult[55]) = "";
		(Bmult[8]  => Cmult[55]) = "";
		(Bmult[9]  => Cmult[55]) = "";
		(Bmult[10] => Cmult[55]) = "";
		(Bmult[11] => Cmult[55]) = "";
		(Bmult[12] => Cmult[55]) = "";
		(Bmult[13] => Cmult[55]) = "";
		(Bmult[14] => Cmult[55]) = "";
		(Bmult[15] => Cmult[55]) = "";
		(Bmult[16] => Cmult[55]) = "";
		(Bmult[17] => Cmult[55]) = "";
		(Bmult[18] => Cmult[55]) = "";
		(Bmult[19] => Cmult[55]) = "";
		(Bmult[20] => Cmult[55]) = "";
		(Bmult[21] => Cmult[55]) = "";
		(Bmult[22] => Cmult[55]) = "";
		(Bmult[23] => Cmult[55]) = "";
		(Bmult[24] => Cmult[55]) = "";
		(Bmult[25] => Cmult[55]) = "";
		(Bmult[26] => Cmult[55]) = "";
		(Bmult[27] => Cmult[55]) = "";
		(Bmult[28] => Cmult[55]) = "";
		(Bmult[29] => Cmult[55]) = "";
		(Bmult[30] => Cmult[55]) = "";
		(Bmult[31] => Cmult[55]) = "";		
		(Valid_mult[0] => Cmult[55]) = "";
		(Valid_mult[1] => Cmult[55]) = "";
		(sel_mul_32x32 => Cmult[55]) = "";
		(Amult[0]  => Cmult[56]) = "";
		(Amult[1]  => Cmult[56]) = "";
		(Amult[2]  => Cmult[56]) = "";
		(Amult[3]  => Cmult[56]) = "";
		(Amult[4]  => Cmult[56]) = "";
		(Amult[5]  => Cmult[56]) = "";
		(Amult[6]  => Cmult[56]) = "";
		(Amult[7]  => Cmult[56]) = "";
		(Amult[8]  => Cmult[56]) = "";
		(Amult[9]  => Cmult[56]) = "";
		(Amult[10] => Cmult[56]) = "";
		(Amult[11] => Cmult[56]) = "";
		(Amult[12] => Cmult[56]) = "";
		(Amult[13] => Cmult[56]) = "";
		(Amult[14] => Cmult[56]) = "";
		(Amult[15] => Cmult[56]) = "";
		(Amult[16] => Cmult[56]) = "";
		(Amult[17] => Cmult[56]) = "";
		(Amult[18] => Cmult[56]) = "";
		(Amult[19] => Cmult[56]) = "";
		(Amult[20] => Cmult[56]) = "";
		(Amult[21] => Cmult[56]) = "";
		(Amult[22] => Cmult[56]) = "";
		(Amult[23] => Cmult[56]) = "";
		(Amult[24] => Cmult[56]) = "";
		(Amult[25] => Cmult[56]) = "";
		(Amult[26] => Cmult[56]) = "";
		(Amult[27] => Cmult[56]) = "";
		(Amult[28] => Cmult[56]) = "";
		(Amult[29] => Cmult[56]) = "";
		(Amult[30] => Cmult[56]) = "";
		(Amult[31] => Cmult[56]) = "";
		(Bmult[0]  => Cmult[56]) = "";
		(Bmult[1]  => Cmult[56]) = "";
		(Bmult[2]  => Cmult[56]) = "";
		(Bmult[3]  => Cmult[56]) = "";
		(Bmult[4]  => Cmult[56]) = "";
		(Bmult[5]  => Cmult[56]) = "";
		(Bmult[6]  => Cmult[56]) = "";
		(Bmult[7]  => Cmult[56]) = "";
		(Bmult[8]  => Cmult[56]) = "";
		(Bmult[9]  => Cmult[56]) = "";
		(Bmult[10] => Cmult[56]) = "";
		(Bmult[11] => Cmult[56]) = "";
		(Bmult[12] => Cmult[56]) = "";
		(Bmult[13] => Cmult[56]) = "";
		(Bmult[14] => Cmult[56]) = "";
		(Bmult[15] => Cmult[56]) = "";
		(Bmult[16] => Cmult[56]) = "";
		(Bmult[17] => Cmult[56]) = "";
		(Bmult[18] => Cmult[56]) = "";
		(Bmult[19] => Cmult[56]) = "";
		(Bmult[20] => Cmult[56]) = "";
		(Bmult[21] => Cmult[56]) = "";
		(Bmult[22] => Cmult[56]) = "";
		(Bmult[23] => Cmult[56]) = "";
		(Bmult[24] => Cmult[56]) = "";
		(Bmult[25] => Cmult[56]) = "";
		(Bmult[26] => Cmult[56]) = "";
		(Bmult[27] => Cmult[56]) = "";
		(Bmult[28] => Cmult[56]) = "";
		(Bmult[29] => Cmult[56]) = "";
		(Bmult[30] => Cmult[56]) = "";
		(Bmult[31] => Cmult[56]) = "";		
		(Valid_mult[0] => Cmult[56]) = "";
		(Valid_mult[1] => Cmult[56]) = "";
		(sel_mul_32x32 => Cmult[56]) = "";
		(Amult[0]  => Cmult[57]) = "";
		(Amult[1]  => Cmult[57]) = "";
		(Amult[2]  => Cmult[57]) = "";
		(Amult[3]  => Cmult[57]) = "";
		(Amult[4]  => Cmult[57]) = "";
		(Amult[5]  => Cmult[57]) = "";
		(Amult[6]  => Cmult[57]) = "";
		(Amult[7]  => Cmult[57]) = "";
		(Amult[8]  => Cmult[57]) = "";
		(Amult[9]  => Cmult[57]) = "";
		(Amult[10] => Cmult[57]) = "";
		(Amult[11] => Cmult[57]) = "";
		(Amult[12] => Cmult[57]) = "";
		(Amult[13] => Cmult[57]) = "";
		(Amult[14] => Cmult[57]) = "";
		(Amult[15] => Cmult[57]) = "";
		(Amult[16] => Cmult[57]) = "";
		(Amult[17] => Cmult[57]) = "";
		(Amult[18] => Cmult[57]) = "";
		(Amult[19] => Cmult[57]) = "";
		(Amult[20] => Cmult[57]) = "";
		(Amult[21] => Cmult[57]) = "";
		(Amult[22] => Cmult[57]) = "";
		(Amult[23] => Cmult[57]) = "";
		(Amult[24] => Cmult[57]) = "";
		(Amult[25] => Cmult[57]) = "";
		(Amult[26] => Cmult[57]) = "";
		(Amult[27] => Cmult[57]) = "";
		(Amult[28] => Cmult[57]) = "";
		(Amult[29] => Cmult[57]) = "";
		(Amult[30] => Cmult[57]) = "";
		(Amult[31] => Cmult[57]) = "";
		(Bmult[0]  => Cmult[57]) = "";
		(Bmult[1]  => Cmult[57]) = "";
		(Bmult[2]  => Cmult[57]) = "";
		(Bmult[3]  => Cmult[57]) = "";
		(Bmult[4]  => Cmult[57]) = "";
		(Bmult[5]  => Cmult[57]) = "";
		(Bmult[6]  => Cmult[57]) = "";
		(Bmult[7]  => Cmult[57]) = "";
		(Bmult[8]  => Cmult[57]) = "";
		(Bmult[9]  => Cmult[57]) = "";
		(Bmult[10] => Cmult[57]) = "";
		(Bmult[11] => Cmult[57]) = "";
		(Bmult[12] => Cmult[57]) = "";
		(Bmult[13] => Cmult[57]) = "";
		(Bmult[14] => Cmult[57]) = "";
		(Bmult[15] => Cmult[57]) = "";
		(Bmult[16] => Cmult[57]) = "";
		(Bmult[17] => Cmult[57]) = "";
		(Bmult[18] => Cmult[57]) = "";
		(Bmult[19] => Cmult[57]) = "";
		(Bmult[20] => Cmult[57]) = "";
		(Bmult[21] => Cmult[57]) = "";
		(Bmult[22] => Cmult[57]) = "";
		(Bmult[23] => Cmult[57]) = "";
		(Bmult[24] => Cmult[57]) = "";
		(Bmult[25] => Cmult[57]) = "";
		(Bmult[26] => Cmult[57]) = "";
		(Bmult[27] => Cmult[57]) = "";
		(Bmult[28] => Cmult[57]) = "";
		(Bmult[29] => Cmult[57]) = "";
		(Bmult[30] => Cmult[57]) = "";
		(Bmult[31] => Cmult[57]) = "";		
		(Valid_mult[0] => Cmult[57]) = "";
		(Valid_mult[1] => Cmult[57]) = "";
		(sel_mul_32x32 => Cmult[57]) = "";
		(Amult[0]  => Cmult[58]) = "";
		(Amult[1]  => Cmult[58]) = "";
		(Amult[2]  => Cmult[58]) = "";
		(Amult[3]  => Cmult[58]) = "";
		(Amult[4]  => Cmult[58]) = "";
		(Amult[5]  => Cmult[58]) = "";
		(Amult[6]  => Cmult[58]) = "";
		(Amult[7]  => Cmult[58]) = "";
		(Amult[8]  => Cmult[58]) = "";
		(Amult[9]  => Cmult[58]) = "";
		(Amult[10] => Cmult[58]) = "";
		(Amult[11] => Cmult[58]) = "";
		(Amult[12] => Cmult[58]) = "";
		(Amult[13] => Cmult[58]) = "";
		(Amult[14] => Cmult[58]) = "";
		(Amult[15] => Cmult[58]) = "";
		(Amult[16] => Cmult[58]) = "";
		(Amult[17] => Cmult[58]) = "";
		(Amult[18] => Cmult[58]) = "";
		(Amult[19] => Cmult[58]) = "";
		(Amult[20] => Cmult[58]) = "";
		(Amult[21] => Cmult[58]) = "";
		(Amult[22] => Cmult[58]) = "";
		(Amult[23] => Cmult[58]) = "";
		(Amult[24] => Cmult[58]) = "";
		(Amult[25] => Cmult[58]) = "";
		(Amult[26] => Cmult[58]) = "";
		(Amult[27] => Cmult[58]) = "";
		(Amult[28] => Cmult[58]) = "";
		(Amult[29] => Cmult[58]) = "";
		(Amult[30] => Cmult[58]) = "";
		(Amult[31] => Cmult[58]) = "";
		(Bmult[0]  => Cmult[58]) = "";
		(Bmult[1]  => Cmult[58]) = "";
		(Bmult[2]  => Cmult[58]) = "";
		(Bmult[3]  => Cmult[58]) = "";
		(Bmult[4]  => Cmult[58]) = "";
		(Bmult[5]  => Cmult[58]) = "";
		(Bmult[6]  => Cmult[58]) = "";
		(Bmult[7]  => Cmult[58]) = "";
		(Bmult[8]  => Cmult[58]) = "";
		(Bmult[9]  => Cmult[58]) = "";
		(Bmult[10] => Cmult[58]) = "";
		(Bmult[11] => Cmult[58]) = "";
		(Bmult[12] => Cmult[58]) = "";
		(Bmult[13] => Cmult[58]) = "";
		(Bmult[14] => Cmult[58]) = "";
		(Bmult[15] => Cmult[58]) = "";
		(Bmult[16] => Cmult[58]) = "";
		(Bmult[17] => Cmult[58]) = "";
		(Bmult[18] => Cmult[58]) = "";
		(Bmult[19] => Cmult[58]) = "";
		(Bmult[20] => Cmult[58]) = "";
		(Bmult[21] => Cmult[58]) = "";
		(Bmult[22] => Cmult[58]) = "";
		(Bmult[23] => Cmult[58]) = "";
		(Bmult[24] => Cmult[58]) = "";
		(Bmult[25] => Cmult[58]) = "";
		(Bmult[26] => Cmult[58]) = "";
		(Bmult[27] => Cmult[58]) = "";
		(Bmult[28] => Cmult[58]) = "";
		(Bmult[29] => Cmult[58]) = "";
		(Bmult[30] => Cmult[58]) = "";
		(Bmult[31] => Cmult[58]) = "";		
		(Valid_mult[0] => Cmult[58]) = "";
		(Valid_mult[1] => Cmult[58]) = "";
		(sel_mul_32x32 => Cmult[58]) = "";	
		(Amult[0]  => Cmult[59]) = "";
		(Amult[1]  => Cmult[59]) = "";
		(Amult[2]  => Cmult[59]) = "";
		(Amult[3]  => Cmult[59]) = "";
		(Amult[4]  => Cmult[59]) = "";
		(Amult[5]  => Cmult[59]) = "";
		(Amult[6]  => Cmult[59]) = "";
		(Amult[7]  => Cmult[59]) = "";
		(Amult[8]  => Cmult[59]) = "";
		(Amult[9]  => Cmult[59]) = "";
		(Amult[10] => Cmult[59]) = "";
		(Amult[11] => Cmult[59]) = "";
		(Amult[12] => Cmult[59]) = "";
		(Amult[13] => Cmult[59]) = "";
		(Amult[14] => Cmult[59]) = "";
		(Amult[15] => Cmult[59]) = "";
		(Amult[16] => Cmult[59]) = "";
		(Amult[17] => Cmult[59]) = "";
		(Amult[18] => Cmult[59]) = "";
		(Amult[19] => Cmult[59]) = "";
		(Amult[20] => Cmult[59]) = "";
		(Amult[21] => Cmult[59]) = "";
		(Amult[22] => Cmult[59]) = "";
		(Amult[23] => Cmult[59]) = "";
		(Amult[24] => Cmult[59]) = "";
		(Amult[25] => Cmult[59]) = "";
		(Amult[26] => Cmult[59]) = "";
		(Amult[27] => Cmult[59]) = "";
		(Amult[28] => Cmult[59]) = "";
		(Amult[29] => Cmult[59]) = "";
		(Amult[30] => Cmult[59]) = "";
		(Amult[31] => Cmult[59]) = "";
		(Bmult[0]  => Cmult[59]) = "";
		(Bmult[1]  => Cmult[59]) = "";
		(Bmult[2]  => Cmult[59]) = "";
		(Bmult[3]  => Cmult[59]) = "";
		(Bmult[4]  => Cmult[59]) = "";
		(Bmult[5]  => Cmult[59]) = "";
		(Bmult[6]  => Cmult[59]) = "";
		(Bmult[7]  => Cmult[59]) = "";
		(Bmult[8]  => Cmult[59]) = "";
		(Bmult[9]  => Cmult[59]) = "";
		(Bmult[10] => Cmult[59]) = "";
		(Bmult[11] => Cmult[59]) = "";
		(Bmult[12] => Cmult[59]) = "";
		(Bmult[13] => Cmult[59]) = "";
		(Bmult[14] => Cmult[59]) = "";
		(Bmult[15] => Cmult[59]) = "";
		(Bmult[16] => Cmult[59]) = "";
		(Bmult[17] => Cmult[59]) = "";
		(Bmult[18] => Cmult[59]) = "";
		(Bmult[19] => Cmult[59]) = "";
		(Bmult[20] => Cmult[59]) = "";
		(Bmult[21] => Cmult[59]) = "";
		(Bmult[22] => Cmult[59]) = "";
		(Bmult[23] => Cmult[59]) = "";
		(Bmult[24] => Cmult[59]) = "";
		(Bmult[25] => Cmult[59]) = "";
		(Bmult[26] => Cmult[59]) = "";
		(Bmult[27] => Cmult[59]) = "";
		(Bmult[28] => Cmult[59]) = "";
		(Bmult[29] => Cmult[59]) = "";
		(Bmult[30] => Cmult[59]) = "";
		(Bmult[31] => Cmult[59]) = "";		
		(Valid_mult[0] => Cmult[59]) = "";
		(Valid_mult[1] => Cmult[59]) = "";
		(sel_mul_32x32 => Cmult[59]) = "";
		(Amult[0]  => Cmult[60]) = "";
		(Amult[1]  => Cmult[60]) = "";
		(Amult[2]  => Cmult[60]) = "";
		(Amult[3]  => Cmult[60]) = "";
		(Amult[4]  => Cmult[60]) = "";
		(Amult[5]  => Cmult[60]) = "";
		(Amult[6]  => Cmult[60]) = "";
		(Amult[7]  => Cmult[60]) = "";
		(Amult[8]  => Cmult[60]) = "";
		(Amult[9]  => Cmult[60]) = "";
		(Amult[10] => Cmult[60]) = "";
		(Amult[11] => Cmult[60]) = "";
		(Amult[12] => Cmult[60]) = "";
		(Amult[13] => Cmult[60]) = "";
		(Amult[14] => Cmult[60]) = "";
		(Amult[15] => Cmult[60]) = "";
		(Amult[16] => Cmult[60]) = "";
		(Amult[17] => Cmult[60]) = "";
		(Amult[18] => Cmult[60]) = "";
		(Amult[19] => Cmult[60]) = "";
		(Amult[20] => Cmult[60]) = "";
		(Amult[21] => Cmult[60]) = "";
		(Amult[22] => Cmult[60]) = "";
		(Amult[23] => Cmult[60]) = "";
		(Amult[24] => Cmult[60]) = "";
		(Amult[25] => Cmult[60]) = "";
		(Amult[26] => Cmult[60]) = "";
		(Amult[27] => Cmult[60]) = "";
		(Amult[28] => Cmult[60]) = "";
		(Amult[29] => Cmult[60]) = "";
		(Amult[30] => Cmult[60]) = "";
		(Amult[31] => Cmult[60]) = "";
		(Bmult[0]  => Cmult[60]) = "";
		(Bmult[1]  => Cmult[60]) = "";
		(Bmult[2]  => Cmult[60]) = "";
		(Bmult[3]  => Cmult[60]) = "";
		(Bmult[4]  => Cmult[60]) = "";
		(Bmult[5]  => Cmult[60]) = "";
		(Bmult[6]  => Cmult[60]) = "";
		(Bmult[7]  => Cmult[60]) = "";
		(Bmult[8]  => Cmult[60]) = "";
		(Bmult[9]  => Cmult[60]) = "";
		(Bmult[10] => Cmult[60]) = "";
		(Bmult[11] => Cmult[60]) = "";
		(Bmult[12] => Cmult[60]) = "";
		(Bmult[13] => Cmult[60]) = "";
		(Bmult[14] => Cmult[60]) = "";
		(Bmult[15] => Cmult[60]) = "";
		(Bmult[16] => Cmult[60]) = "";
		(Bmult[17] => Cmult[60]) = "";
		(Bmult[18] => Cmult[60]) = "";
		(Bmult[19] => Cmult[60]) = "";
		(Bmult[20] => Cmult[60]) = "";
		(Bmult[21] => Cmult[60]) = "";
		(Bmult[22] => Cmult[60]) = "";
		(Bmult[23] => Cmult[60]) = "";
		(Bmult[24] => Cmult[60]) = "";
		(Bmult[25] => Cmult[60]) = "";
		(Bmult[26] => Cmult[60]) = "";
		(Bmult[27] => Cmult[60]) = "";
		(Bmult[28] => Cmult[60]) = "";
		(Bmult[29] => Cmult[60]) = "";
		(Bmult[30] => Cmult[60]) = "";
		(Bmult[31] => Cmult[60]) = "";		
		(Valid_mult[0] => Cmult[60]) = "";
		(Valid_mult[1] => Cmult[60]) = "";
		(sel_mul_32x32 => Cmult[60]) = "";
		(Amult[0]  => Cmult[61]) = "";
		(Amult[1]  => Cmult[61]) = "";
		(Amult[2]  => Cmult[61]) = "";
		(Amult[3]  => Cmult[61]) = "";
		(Amult[4]  => Cmult[61]) = "";
		(Amult[5]  => Cmult[61]) = "";
		(Amult[6]  => Cmult[61]) = "";
		(Amult[7]  => Cmult[61]) = "";
		(Amult[8]  => Cmult[61]) = "";
		(Amult[9]  => Cmult[61]) = "";
		(Amult[10] => Cmult[61]) = "";
		(Amult[11] => Cmult[61]) = "";
		(Amult[12] => Cmult[61]) = "";
		(Amult[13] => Cmult[61]) = "";
		(Amult[14] => Cmult[61]) = "";
		(Amult[15] => Cmult[61]) = "";
		(Amult[16] => Cmult[61]) = "";
		(Amult[17] => Cmult[61]) = "";
		(Amult[18] => Cmult[61]) = "";
		(Amult[19] => Cmult[61]) = "";
		(Amult[20] => Cmult[61]) = "";
		(Amult[21] => Cmult[61]) = "";
		(Amult[22] => Cmult[61]) = "";
		(Amult[23] => Cmult[61]) = "";
		(Amult[24] => Cmult[61]) = "";
		(Amult[25] => Cmult[61]) = "";
		(Amult[26] => Cmult[61]) = "";
		(Amult[27] => Cmult[61]) = "";
		(Amult[28] => Cmult[61]) = "";
		(Amult[29] => Cmult[61]) = "";
		(Amult[30] => Cmult[61]) = "";
		(Amult[31] => Cmult[61]) = "";
		(Bmult[0]  => Cmult[61]) = "";
		(Bmult[1]  => Cmult[61]) = "";
		(Bmult[2]  => Cmult[61]) = "";
		(Bmult[3]  => Cmult[61]) = "";
		(Bmult[4]  => Cmult[61]) = "";
		(Bmult[5]  => Cmult[61]) = "";
		(Bmult[6]  => Cmult[61]) = "";
		(Bmult[7]  => Cmult[61]) = "";
		(Bmult[8]  => Cmult[61]) = "";
		(Bmult[9]  => Cmult[61]) = "";
		(Bmult[10] => Cmult[61]) = "";
		(Bmult[11] => Cmult[61]) = "";
		(Bmult[12] => Cmult[61]) = "";
		(Bmult[13] => Cmult[61]) = "";
		(Bmult[14] => Cmult[61]) = "";
		(Bmult[15] => Cmult[61]) = "";
		(Bmult[16] => Cmult[61]) = "";
		(Bmult[17] => Cmult[61]) = "";
		(Bmult[18] => Cmult[61]) = "";
		(Bmult[19] => Cmult[61]) = "";
		(Bmult[20] => Cmult[61]) = "";
		(Bmult[21] => Cmult[61]) = "";
		(Bmult[22] => Cmult[61]) = "";
		(Bmult[23] => Cmult[61]) = "";
		(Bmult[24] => Cmult[61]) = "";
		(Bmult[25] => Cmult[61]) = "";
		(Bmult[26] => Cmult[61]) = "";
		(Bmult[27] => Cmult[61]) = "";
		(Bmult[28] => Cmult[61]) = "";
		(Bmult[29] => Cmult[61]) = "";
		(Bmult[30] => Cmult[61]) = "";
		(Bmult[31] => Cmult[61]) = "";		
		(Valid_mult[0] => Cmult[61]) = "";
		(Valid_mult[1] => Cmult[61]) = "";
		(sel_mul_32x32 => Cmult[61]) = "";
		(Amult[0]  => Cmult[62]) = "";
		(Amult[1]  => Cmult[62]) = "";
		(Amult[2]  => Cmult[62]) = "";
		(Amult[3]  => Cmult[62]) = "";
		(Amult[4]  => Cmult[62]) = "";
		(Amult[5]  => Cmult[62]) = "";
		(Amult[6]  => Cmult[62]) = "";
		(Amult[7]  => Cmult[62]) = "";
		(Amult[8]  => Cmult[62]) = "";
		(Amult[9]  => Cmult[62]) = "";
		(Amult[10] => Cmult[62]) = "";
		(Amult[11] => Cmult[62]) = "";
		(Amult[12] => Cmult[62]) = "";
		(Amult[13] => Cmult[62]) = "";
		(Amult[14] => Cmult[62]) = "";
		(Amult[15] => Cmult[62]) = "";
		(Amult[16] => Cmult[62]) = "";
		(Amult[17] => Cmult[62]) = "";
		(Amult[18] => Cmult[62]) = "";
		(Amult[19] => Cmult[62]) = "";
		(Amult[20] => Cmult[62]) = "";
		(Amult[21] => Cmult[62]) = "";
		(Amult[22] => Cmult[62]) = "";
		(Amult[23] => Cmult[62]) = "";
		(Amult[24] => Cmult[62]) = "";
		(Amult[25] => Cmult[62]) = "";
		(Amult[26] => Cmult[62]) = "";
		(Amult[27] => Cmult[62]) = "";
		(Amult[28] => Cmult[62]) = "";
		(Amult[29] => Cmult[62]) = "";
		(Amult[30] => Cmult[62]) = "";
		(Amult[31] => Cmult[62]) = "";
		(Bmult[0]  => Cmult[62]) = "";
		(Bmult[1]  => Cmult[62]) = "";
		(Bmult[2]  => Cmult[62]) = "";
		(Bmult[3]  => Cmult[62]) = "";
		(Bmult[4]  => Cmult[62]) = "";
		(Bmult[5]  => Cmult[62]) = "";
		(Bmult[6]  => Cmult[62]) = "";
		(Bmult[7]  => Cmult[62]) = "";
		(Bmult[8]  => Cmult[62]) = "";
		(Bmult[9]  => Cmult[62]) = "";
		(Bmult[10] => Cmult[62]) = "";
		(Bmult[11] => Cmult[62]) = "";
		(Bmult[12] => Cmult[62]) = "";
		(Bmult[13] => Cmult[62]) = "";
		(Bmult[14] => Cmult[62]) = "";
		(Bmult[15] => Cmult[62]) = "";
		(Bmult[16] => Cmult[62]) = "";
		(Bmult[17] => Cmult[62]) = "";
		(Bmult[18] => Cmult[62]) = "";
		(Bmult[19] => Cmult[62]) = "";
		(Bmult[20] => Cmult[62]) = "";
		(Bmult[21] => Cmult[62]) = "";
		(Bmult[22] => Cmult[62]) = "";
		(Bmult[23] => Cmult[62]) = "";
		(Bmult[24] => Cmult[62]) = "";
		(Bmult[25] => Cmult[62]) = "";
		(Bmult[26] => Cmult[62]) = "";
		(Bmult[27] => Cmult[62]) = "";
		(Bmult[28] => Cmult[62]) = "";
		(Bmult[29] => Cmult[62]) = "";
		(Bmult[30] => Cmult[62]) = "";
		(Bmult[31] => Cmult[62]) = "";		
		(Valid_mult[0] => Cmult[62]) = "";
		(Valid_mult[1] => Cmult[62]) = "";
		(sel_mul_32x32 => Cmult[62]) = "";
		(Amult[0]  => Cmult[63]) = "";
		(Amult[1]  => Cmult[63]) = "";
		(Amult[2]  => Cmult[63]) = "";
		(Amult[3]  => Cmult[63]) = "";
		(Amult[4]  => Cmult[63]) = "";
		(Amult[5]  => Cmult[63]) = "";
		(Amult[6]  => Cmult[63]) = "";
		(Amult[7]  => Cmult[63]) = "";
		(Amult[8]  => Cmult[63]) = "";
		(Amult[9]  => Cmult[63]) = "";
		(Amult[10] => Cmult[63]) = "";
		(Amult[11] => Cmult[63]) = "";
		(Amult[12] => Cmult[63]) = "";
		(Amult[13] => Cmult[63]) = "";
		(Amult[14] => Cmult[63]) = "";
		(Amult[15] => Cmult[63]) = "";
		(Amult[16] => Cmult[63]) = "";
		(Amult[17] => Cmult[63]) = "";
		(Amult[18] => Cmult[63]) = "";
		(Amult[19] => Cmult[63]) = "";
		(Amult[20] => Cmult[63]) = "";
		(Amult[21] => Cmult[63]) = "";
		(Amult[22] => Cmult[63]) = "";
		(Amult[23] => Cmult[63]) = "";
		(Amult[24] => Cmult[63]) = "";
		(Amult[25] => Cmult[63]) = "";
		(Amult[26] => Cmult[63]) = "";
		(Amult[27] => Cmult[63]) = "";
		(Amult[28] => Cmult[63]) = "";
		(Amult[29] => Cmult[63]) = "";
		(Amult[30] => Cmult[63]) = "";
		(Amult[31] => Cmult[63]) = "";
		(Bmult[0]  => Cmult[63]) = "";
		(Bmult[1]  => Cmult[63]) = "";
		(Bmult[2]  => Cmult[63]) = "";
		(Bmult[3]  => Cmult[63]) = "";
		(Bmult[4]  => Cmult[63]) = "";
		(Bmult[5]  => Cmult[63]) = "";
		(Bmult[6]  => Cmult[63]) = "";
		(Bmult[7]  => Cmult[63]) = "";
		(Bmult[8]  => Cmult[63]) = "";
		(Bmult[9]  => Cmult[63]) = "";
		(Bmult[10] => Cmult[63]) = "";
		(Bmult[11] => Cmult[63]) = "";
		(Bmult[12] => Cmult[63]) = "";
		(Bmult[13] => Cmult[63]) = "";
		(Bmult[14] => Cmult[63]) = "";
		(Bmult[15] => Cmult[63]) = "";
		(Bmult[16] => Cmult[63]) = "";
		(Bmult[17] => Cmult[63]) = "";
		(Bmult[18] => Cmult[63]) = "";
		(Bmult[19] => Cmult[63]) = "";
		(Bmult[20] => Cmult[63]) = "";
		(Bmult[21] => Cmult[63]) = "";
		(Bmult[22] => Cmult[63]) = "";
		(Bmult[23] => Cmult[63]) = "";
		(Bmult[24] => Cmult[63]) = "";
		(Bmult[25] => Cmult[63]) = "";
		(Bmult[26] => Cmult[63]) = "";
		(Bmult[27] => Cmult[63]) = "";
		(Bmult[28] => Cmult[63]) = "";
		(Bmult[29] => Cmult[63]) = "";
		(Bmult[30] => Cmult[63]) = "";
		(Bmult[31] => Cmult[63]) = "";		
		(Valid_mult[0] => Cmult[63]) = "";
		(Valid_mult[1] => Cmult[63]) = "";
		(sel_mul_32x32 => Cmult[63]) = "";		
    endspecify
`endif
	
	always @(*) begin
		if (sel_mul_32x32 == 1'b1) begin
			if (Valid_mult[0] == 1'b1) begin
				Cmult <= Amult * Bmult;
			end
		end else begin
			if (Valid_mult[0] == 1'b1) begin
				Cmult[31:0] <= Amult[15:0] * Bmult[15:0];
			end
			if (Valid_mult[1] == 1'b1) begin
				Cmult[63:32] <= Amult[31:16] * Bmult[31:16];
			end
		end
	end


endmodule
