(* blackbox *)
module CYINIT_CONSTANTS(
	C0, C1
);
	output wire C0;
	output wire C1;

  assign C0 = 0;
  assign C1 = 1;
endmodule

