module top(input i0, input i1, input i2, output o0, output o1, output o2, output o3, output o4, output o5);
   assign o0 = i0;
   assign o1 = i1;
   assign o2 = i1;
   assign o3 = i2;
   assign o4 = i2;
   assign o5 = i2;
endmodule // top
