(* whitebox *)
module TIEOFF(
	HARD0, HARD1
);
	output wire HARD0;
	output wire HARD1;

  assign HARD0 = 0;
  assign HARD1 = 1;
endmodule
