module top(
    input  wire clk,

    output [3:0] wire led
);
  assign led = 4'b1010;
endmodule
