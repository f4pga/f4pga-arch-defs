module data_generator(
    input  wire CLK,
    input  wire CE,
    output wire D1,
    output wire D2
);

    // Ring buffers
    reg [254:0] ring1;
    initial ring1 <= 255'b010100110101100010111100101101010010011100001110110010000001011011011111011000101110100111001101101100110111101100001111100110000001011011010000111011000010001010101000101111101110110111100110110000001100101111111011010111100001101100001101111111001110111;

    reg [255:0] ring2;
    initial ring2 <= 256'b1010101100101110000100100101010000100000101110111011110111011111000111101101010101110111010011011101100100011111111101101000111110110110100010011011001001000011100011001001110001110101000001010011011001100101000001011111011101010000110011101111110100110010;

    reg [256:0] ring3;
    initial ring3 <= 257'b10000001100111000110101001001111100011011001100011011111000100110100110001011101100111110101101111101011000101110100100110110010000111100011111101010000000100101000100100110101011111011000100100001001100110101011111101101011011100010101000111110010110011110;

    // Rotate ring buffers
    always @(posedge CLK)
        if (CE) ring1 <= {ring1[0], ring1[254:1]};
    always @(posedge CLK)
        if (CE) ring2 <= {ring2[0], ring2[255:1]};
    always @(posedge CLK)
        if (CE) ring3 <= {ring3[0], ring3[256:1]};

    // Output data
    assign D1 = ring1[0] ^ ring2[0];
    assign D2 = ring2[0] ^ ring3[0];

endmodule
