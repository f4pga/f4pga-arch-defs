`timescale 1ns/10ps
(* blackbox *)
(* keep *)
module ASSPL (
  input  wire        SEL_18_top,
  input  wire        SEL_18_bottom,
  input  wire        SEL_18_left,
  input  wire        SEL_18_right,
  input  wire        SPI_CLK,
  input  wire        default_SPI_IO_mux,
  input  wire        SPI_SSn,
  input  wire        SPI_MOSI,
  input  wire        RAM8K_P1_mux,
  input  wire [3:0]  RAM8K_RM_af,
  input  wire        RAM8K_RME_af,
  input  wire        RAM8K_P0_CLK,
  input  wire [3:0]  af_burnin_mode,
  input  wire        osc_en,
  input  wire        osc_fsel,
  input  wire [2:0]  osc_sel,
  input  wire [16:0] RAM8K_P0_WR_DATA,
  input  wire [1:0]  RAM8K_P0_WR_BE,
  input  wire        af_spi_cpha,
  input  wire        af_spi_cpol,
  input  wire        af_spi_lsbf,
  input  wire        RAM8K_P0_WR_EN,
  input  wire        RAM8K_TEST1_af,
  input  wire [11:0] RAM8K_P0_ADDR,
  input  wire        RAM8K_P1_CLK,
  input  wire [11:0] RAM8K_P1_ADDR,
  input  wire        RAM8K_P1_RD_EN,
  input  wire        RESET_n,
  input  wire        RAM8K_fifo_en,
  input  wire [7:0]  int_i,
  input  wire        reg_clk_int,
  input  wire        reg_wr_en_int,
  input  wire        reg_rd_en_int,
  input  wire [7:0]  reg_wr_data_int,
  input  wire        drive_io_en_4,
  input  wire        drive_io_en_5,
  input  wire [1:0]  reg_addr_int,
  input  wire [6:0]  A2F_Status,
  input  wire        af_fpga_int_en,
  input  wire [31:0] af_dev_id,
  input  wire [7:0]  A2F_GP_IN,
  input  wire [7:0]  A2F_RD_DATA,
  input  wire        A2F_ACK,
  input  wire [31:0] Amult0,
  input  wire        drive_io_en_2,
  input  wire        drive_io_en_3,
  input  wire        drive_io_en_0,
  input  wire        drive_io_en_1,
  input  wire [31:0] Bmult0,
  input  wire        RAM0_CLK,
  input  wire        Valid_mult0,
  input  wire        af_opt_0,
  input  wire        af_opt_1,
  input  wire [3:0]  RAM0_RM_af,
  input  wire        RAM0_RME_af,
  input  wire        \af_plat_id[0] ,
  input  wire        \af_plat_id[1] ,
  input  wire        \af_plat_id[2] ,
  input  wire        \af_plat_id[3] ,
  input  wire        \af_plat_id[4] ,
  input  wire        \af_plat_id[5] ,
  input  wire        \af_plat_id[6] ,
  input  wire        \af_plat_id[7] ,
  input  wire [35:0] RAM0_WR_DATA,
  input  wire [3:0]  RAM0_WR_BE,
  input  wire        RAM0_RD_EN,
  input  wire        RAM0_WR_EN,
  input  wire        RAM0_TEST1_af,
  input  wire [8:0]  RAM0_ADDR,
  output wire        SPI_MISO,
  output wire        SPI_MISOe,
  output wire [16:0] RAM8K_P1_RD_DATA,
  output wire        SYSCLK_x2,
  output wire        SYSCLK,
  output wire        fast_clk_out,
  output wire        RAM8K_fifo_almost_full,
  output wire [3:0]  RAM8K_fifo_full_flag,
  output wire        RAM8K_fifo_almost_empty,
  output wire [3:0]  RAM8K_fifo_empty_flag,
  output wire        int_o,
  output wire [7:0]  reg_rd_data_int,
  output wire [7:0]  A2F_Control,
  output wire [7:0]  A2F_GP_OUT,
  output wire        A2F_REQ,
  output wire        A2F_RWn,
  output wire [7:0]  A2F_WR_DATA,
  output wire [7:0]  A2F_ADDR,
  output wire [63:0] Cmult0,
  output wire [35:0] RAM0_RD_DATA
);

endmodule
