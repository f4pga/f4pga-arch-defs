module IBUF (
  input  I,
  output O
);

  assign O = I;

endmodule


module OBUF (
  input  I,
  output O
);

  assign O = I;

endmodule

