(* whitebox *)
(* MODEL_NAME="logic_0" *)
module LOGIC_0_CELL (
    output wire a
);

    assign a = 1'b0;

endmodule
