(* whitebox *)
module FDPE(D, SR, CE, CLK, Q);
    input  D;
    input  SR;
    input  CE;
    input  CLK;
    output  Q;
endmodule
