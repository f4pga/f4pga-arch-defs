`ifdef af512x16_512x16
`else
`define af512x16_512x16
/************************************************************************
** File : af512x16_512x16.v
** Design Date: April 11, 2005
** Creation Date: Thu Dec 06 23:09:33 2012

** Created By SpDE Version: SpDE 2012.1.1 Release Build
** Author: QuickLogic India Development Centre,
** Copyright (C) 1998, Customers of QuickLogic may copy and modify this
** file for use in designing QuickLogic devices only.
** Description : This file is autogenerated RTL code that describes the
** top level design file for Asynchronous FIFO using QuickLogic's
** RAM block resources.
************************************************************************/
module af512x16_512x16(DIN,Fifo_Push_Flush,Fifo_Pop_Flush,PUSH,POP,Push_Clk,Pop_Clk,
       Push_Clk_En,Pop_Clk_En,Push_Clk_Sel,Pop_Clk_Sel,Fifo_Dir,Async_Flush,Async_Flush_Sel,
       Almost_Full,Almost_Empty,PUSH_FLAG,POP_FLAG,DOUT);


input Fifo_Push_Flush,Fifo_Pop_Flush;
input Push_Clk,Pop_Clk;
input PUSH,POP;
input [15:0] DIN;
input Push_Clk_En,Pop_Clk_En,Push_Clk_Sel,Pop_Clk_Sel,Fifo_Dir,Async_Flush,Async_Flush_Sel;
output [15:0] DOUT;
output [3:0] PUSH_FLAG,POP_FLAG;
output Almost_Full,Almost_Empty;

parameter wr_depth_int = 512;
parameter rd_depth_int = 512;
parameter wr_width_int = 16;
parameter rd_width_int = 16;
parameter reg_rd_int = 0;
parameter sync_fifo_int = 0;

supply0 GND;
supply1 VCC;

assign DOUT = DIN;
assign PUSH_FLAG = {Fifo_Push_Flush,Fifo_Pop_Flush,Push_Clk,Pop_Clk};
assign POP_FLAG = {Push_Clk_En,Pop_Clk_En,Push_Clk_Sel,Pop_Clk_Sel};
assign Almost_Full = Fifo_Dir;
assign Almost_Empty = Async_Flush_Sel;

endmodule
`endif
