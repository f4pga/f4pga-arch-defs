(* whitebox *)
module FF(D, SR, CE, CLK, Q);
    input D;
    input SR;
    input CE;
    input CLK;
    output Q;
endmodule
