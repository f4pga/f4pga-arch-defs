`timescale 1ps/1ps
(* whitebox *)
module GND (
    output wire GND
);

    assign GND = 1'b0;

endmodule
