(* CLASS="input" *)
module VPR_IPAD(inpad);
    output wire inpad;

endmodule
