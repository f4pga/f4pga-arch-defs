module  \$_DFF_N_ (input D, C, output Q); FF _TECHMAP_REPLACE_ (.D(D), .Q(Q), .clk(C)); endmodule
module  \$_DFF_P_ (input D, C, output Q); FF _TECHMAP_REPLACE_ (.D(D), .Q(Q), .clk(C)); endmodule
