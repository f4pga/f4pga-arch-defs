(* whitebox *)
module CE_VCC(CE_OUT);
    output wire CE_OUT;

    assign CE_OUT = 1;
endmodule
