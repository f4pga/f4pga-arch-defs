module top(
	input [11:0] in,
	output [11:0] out
);

assign out = in;

endmodule
