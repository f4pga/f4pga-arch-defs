(* whitebox *)
module SR_USED(SR, SR_OUT);
    input wire SR;
    output wire SR_OUT;

    assign SR_OUT = SR;
endmodule
