(* CLASS="lut" *)
(* whitebox *)
module LUT5 (in, out);
    (* PORT_CLASS="lut_in" *)
    input wire [4:0] in;
    (* PORT_CLASS="lut_out" *)
    output wire out;
endmodule
