(* whitebox *)
(* MODEL_NAME="logic_1" *)
module LOGIC_1_CELL (
    output wire a
);

    assign a = 1'b1;

endmodule
