module top(
	output wire [3:0] led,
	input wire rx,
	output wire tx,
	input wire clk125
);

	wire [3:0] fclk;
	wire [3:0] fresetn;
	wire reset;
	wire [1:0] gpios;
	wire [19:0] irqf2p;
	wire fclk0_bg;

	/* Master AXI bus */
	/* AR */
	wire [31:0] MAXIGP0ARADDR;
	wire MAXIGP0ARCACHE;
	wire MAXIGP0ARVALID;
	wire [2:0] MAXIGP0ARPROT;
	wire MAXIGP0ARREADY;
	wire [11:0] MAXIGP0ARID;
	/* AW */
	wire [31:0] MAXIGP0AWADDR;
	wire MAXIGP0AWVALID;
	wire [2:0] MAXIGP0AWPROT;
	wire MAXIGP0AWREADY;
	wire [11:0] MAXIGP0AWID;
	/* B */
	wire MAXIGP0BREADY;
	wire [1:0] MAXIGP0BRESP;
	wire MAXIGP0BVALID;
	wire [11:0] MAXIGP0BID;
	/* W */
	wire MAXIGP0RREADY;
	wire [31:0] MAXIGP0WDATA;
	wire [3:0] MAXIGP0WSTRB;
	wire MAXIGP0WVALID;
	wire MAXIGP0WREADY;
	wire [11:0] MAXIGP0WID;
	/* R */
	wire [31:0] MAXIGP0RDATA;
	wire [1:0] MAXIGP0RRESP;
	wire MAXIGP0RVALID;
	wire [11:0] MAXIGP0RID;

	/* PS7 Inputs */
	wire MAXIGP0ACLK;

	/* Slave AXI bus */
	wire SAXIGP0ACLK;
	wire MAXIGP0ARESETN;

	/* AR */
	wire [31:0] SAXIGP0ARADDR;
	wire [1:0]  SAXIGP0ARBURST;
	wire [3:0]  SAXIGP0ARCACHE;
	wire [11:0] SAXIGP0ARID;
	wire [3:0]  SAXIGP0ARLEN;
	wire [1:0]  SAXIGP0ARLOCK;
	wire [2:0]  SAXIGP0ARPROT;
	wire [3:0]  SAXIGP0ARQOS;
	wire [1:0]  SAXIGP0ARSIZE;
	wire SAXIGP0ARVALID;
	wire SAXIGP0ARREADY;
	/* AW */
	wire [31:0] SAXIGP0AWADDR;
	wire [1:0]  SAXIGP0AWBURST;
	wire [3:0]  SAXIGP0AWCACHE;
	wire [11:0] SAXIGP0AWID;
	wire [3:0]  SAXIGP0AWLEN;
	wire [1:0]  SAXIGP0AWLOCK;
	wire [2:0]  SAXIGP0AWPROT;
	wire [3:0]  SAXIGP0AWQOS;
	wire [1:0]  SAXIGP0AWSIZE;
	wire SAXIGP0AWVALID;
	wire SAXIGP0AWREADY;
	/* B */
	wire [11:0] SAXIGP0BID;
	wire [1:0]  SAXIGP0BRESP;
	wire SAXIGP0BVALID;
	wire SAXIGP0BREADY;
	/* R */
	wire [31:0] SAXIGP0RDATA;
	wire [11:0] SAXIGP0RID;
	wire [1:0] SAXIGP0RRESP;
	wire SAXIGP0RLAST;
	wire SAXIGP0RVALID;
	wire SAXIGP0RREADY;
	/* W */
	wire [31:0] SAXIGP0WDATA;
	wire [11:0] SAXIGP0WID;
	wire [3:0]  SAXIGP0WSTRB;
	wire SAXIGP0WVALID;
	wire SAXIGP0WLAST;
	wire SAXIGP0WREADY;

	wire litex_reset;

	assign reset_maxi_gp0 = ~fresetn[0];
	assign litex_reset = ~(SAXIGP0ARESETN & gpios[0]);
	assign SAXIGP0ACLK = fclk0_bg;
	assign MAXIGP0ACLK = fclk0_bg;
	assign irqf2p = 20'h00000;

	reg [31:0] counter;

	always @(posedge fclk0_bg)
	if(reset) begin
		counter <= 32'h00000000;
	end else begin
		counter <= counter + 1'b1;
		if(counter == 32'hffffffff) begin
			counter <= 32'h00000000;
		end
	end

	assign led[0] = gpios[0];
	assign led[1] = litex_reset;
	assign led[2] = reset;
	assign led[3] = counter[23];

    BUFG bg (
	.I(clk125),
	.O(clk125_bg)
    );

    // The PS7
    (* KEEP, DONT_TOUCH *)
    PS7 the_PS (
	.DMA0DATYPE			(),
	.DMA0DAVALID			(),
	.DMA0DRREADY			(),
	.DMA0RSTN			(),
	.DMA1DATYPE			(),
	.DMA1DAVALID			(),
	.DMA1DRREADY			(),
	.DMA1RSTN			(),
	.DMA2DATYPE			(),
	.DMA2DAVALID			(),
	.DMA2DRREADY			(),
	.DMA2RSTN			(),
	.DMA3DATYPE			(),
	.DMA3DAVALID			(),
	.DMA3DRREADY			(),
	.DMA3RSTN			(),
	.EMIOCAN0PHYTX			(),
	.EMIOCAN1PHYTX			(),
	.EMIOENET0GMIITXD		(),
	.EMIOENET0GMIITXEN		(),
	.EMIOENET0GMIITXER		(),
	.EMIOENET0MDIOMDC		(),
	.EMIOENET0MDIOO			(),
	.EMIOENET0MDIOTN		(),
	.EMIOENET0PTPDELAYREQRX		(),
	.EMIOENET0PTPDELAYREQTX		(),
	.EMIOENET0PTPPDELAYREQRX	(),
	.EMIOENET0PTPPDELAYREQTX	(),
	.EMIOENET0PTPPDELAYRESPRX	(),
	.EMIOENET0PTPPDELAYRESPTX	(),
	.EMIOENET0PTPSYNCFRAMERX	(),
	.EMIOENET0PTPSYNCFRAMETX	(),
	.EMIOENET0SOFRX			(),
	.EMIOENET0SOFTX			(),
	.EMIOENET1GMIITXD		(),
	.EMIOENET1GMIITXEN		(),
	.EMIOENET1GMIITXER		(),
	.EMIOENET1MDIOMDC		(),
	.EMIOENET1MDIOO			(),
	.EMIOENET1MDIOTN		(),
	.EMIOENET1PTPDELAYREQRX		(),
	.EMIOENET1PTPDELAYREQTX		(),
	.EMIOENET1PTPPDELAYREQRX	(),
	.EMIOENET1PTPPDELAYREQTX	(),
	.EMIOENET1PTPPDELAYRESPRX	(),
	.EMIOENET1PTPPDELAYRESPTX	(),
	.EMIOENET1PTPSYNCFRAMERX	(),
	.EMIOENET1PTPSYNCFRAMETX	(),
	.EMIOENET1SOFRX			(),
	.EMIOENET1SOFTX			(),
	.EMIOGPIOO			(),
	.EMIOGPIOTN			(),
	.EMIOI2C0SCLO			(),
	.EMIOI2C0SCLTN			(),
	.EMIOI2C0SDAO			(),
	.EMIOI2C0SDATN			(),
	.EMIOI2C1SCLO			(),
	.EMIOI2C1SCLTN			(),
	.EMIOI2C1SDAO			(),
	.EMIOI2C1SDATN			(),
	.EMIOPJTAGTDO			(),
	.EMIOPJTAGTDTN			(),
	.EMIOSDIO0BUSPOW		(),
	.EMIOSDIO0BUSVOLT		(),
	.EMIOSDIO0CLK			(),
	.EMIOSDIO0CMDO			(),
	.EMIOSDIO0CMDTN			(),
	.EMIOSDIO0DATAO			(),
	.EMIOSDIO0DATATN		(),
	.EMIOSDIO0LED			(),
	.EMIOSDIO1BUSPOW		(),
	.EMIOSDIO1BUSVOLT		(),
	.EMIOSDIO1CLK			(),
	.EMIOSDIO1CMDO			(),
	.EMIOSDIO1CMDTN			(),
	.EMIOSDIO1DATAO			(),
	.EMIOSDIO1DATATN		(),
	.EMIOSDIO1LED			(),
	.EMIOSPI0MO			(),
	.EMIOSPI0MOTN			(),
	.EMIOSPI0SCLKO			(),
	.EMIOSPI0SCLKTN			(),
	.EMIOSPI0SO		   (),
	.EMIOSPI0SSNTN			(),
	.EMIOSPI0SSON			(),
	.EMIOSPI0STN			(),
	.EMIOSPI1MO			    (),
	.EMIOSPI1MOTN			(),
	.EMIOSPI1SCLKO			(),
	.EMIOSPI1SCLKTN			(),
	.EMIOSPI1SO			    (),
	.EMIOSPI1SSNTN			(),
	.EMIOSPI1SSON			(),
	.EMIOSPI1STN			(),
	.EMIOTRACECTL			(),
	.EMIOTRACEDATA			(),
	.EMIOTTC0WAVEO			(),
	.EMIOTTC1WAVEO			(),
	.EMIOUART0DTRN			(),
	.EMIOUART0RTSN			(),
	.EMIOUART0TX			(),
	.EMIOUART1DTRN			(),
	.EMIOUART1RTSN			(),
	.EMIOUART1TX			(),
	.EMIOUSB0PORTINDCTL		(),
	.EMIOUSB0VBUSPWRSELECT	(),
	.EMIOUSB1PORTINDCTL		(),
	.EMIOUSB1VBUSPWRSELECT	(),
	.EMIOWDTRSTO			(),
	.EVENTEVENTO			(),
	.EVENTSTANDBYWFE		(),
	.EVENTSTANDBYWFI		(),
	.FCLKCLK			    (fclk),
	.FCLKRESETN			    (fresetn),
	.FTMTF2PTRIGACK			(),
	.FTMTP2FDEBUG			(),
	.FTMTP2FTRIG			(),
	.IRQP2F				(),
	.MAXIGP0ARADDR			(MAXIGP0ARADDR	),
	.MAXIGP0ARBURST			(),
	.MAXIGP0ARCACHE			(),
	.MAXIGP0ARESETN			(),
	.MAXIGP0ARID			(MAXIGP0ARID),
	.MAXIGP0ARLEN			(),
	.MAXIGP0ARLOCK			(),
	.MAXIGP0ARPROT			(MAXIGP0ARPROT	),
	.MAXIGP0ARQOS			(),
	.MAXIGP0ARSIZE			(),
	.MAXIGP0ARVALID			(MAXIGP0ARVALID	),
	.MAXIGP0AWADDR			(MAXIGP0AWADDR	),
	.MAXIGP0AWBURST			(),
	.MAXIGP0AWCACHE			(),
	.MAXIGP0AWID			(MAXIGP0AWID),
	.MAXIGP0AWLEN			(),
	.MAXIGP0AWLOCK			(),
	.MAXIGP0AWPROT			(MAXIGP0AWPROT),
	.MAXIGP0AWQOS			(),
	.MAXIGP0AWSIZE			(),
	.MAXIGP0AWVALID			(MAXIGP0AWVALID	),
	.MAXIGP0BREADY			(MAXIGP0BREADY	),
	.MAXIGP0RREADY			(MAXIGP0RREADY	),
	.MAXIGP0WDATA			(MAXIGP0WDATA	),
	.MAXIGP0WID			(MAXIGP0WID),
	.MAXIGP0WLAST			(),
	.MAXIGP0WSTRB			(MAXIGP0WSTRB	),
	.MAXIGP0WVALID			(MAXIGP0WVALID	),
	.MAXIGP1ARADDR			(),
	.MAXIGP1ARBURST			(),
	.MAXIGP1ARCACHE			(),
	.MAXIGP1ARESETN			(),
	.MAXIGP1ARID			(),
	.MAXIGP1ARLEN			(),
	.MAXIGP1ARLOCK			(),
	.MAXIGP1ARPROT			(),
	.MAXIGP1ARQOS			(),
	.MAXIGP1ARSIZE			(),
	.MAXIGP1ARVALID			(),
	.MAXIGP1AWADDR			(),
	.MAXIGP1AWBURST			(),
	.MAXIGP1AWCACHE			(),
	.MAXIGP1AWID			(),
	.MAXIGP1AWLEN			(),
	.MAXIGP1AWLOCK			(),
	.MAXIGP1AWPROT			(),
	.MAXIGP1AWQOS			(),
	.MAXIGP1AWSIZE			(),
	.MAXIGP1AWVALID			(),
	.MAXIGP1BREADY			(),
	.MAXIGP1RREADY			(),
	.MAXIGP1WDATA			(),
	.MAXIGP1WID			(),
	.MAXIGP1WLAST			(),
	.MAXIGP1WSTRB			(),
	.MAXIGP1WVALID			(),
	.SAXIACPARESETN			(),
	.SAXIACPARREADY			(),
	.SAXIACPAWREADY			(),
	.SAXIACPBID			(),
	.SAXIACPBRESP			(),
	.SAXIACPBVALID			(),
	.SAXIACPRDATA			(),
	.SAXIACPRID			(),
	.SAXIACPRLAST			(),
	.SAXIACPRRESP			(),
	.SAXIACPRVALID			(),
	.SAXIACPWREADY			(),
	/* SAXI GP0 outputs */
	.SAXIGP1ARESETN			(SAXIGP0ARESETN ),
	.SAXIGP1ARREADY			(SAXIGP0ARREADY	),
	.SAXIGP1AWREADY			(SAXIGP0AWREADY	),
	.SAXIGP1BID			(SAXIGP0BID	),
	.SAXIGP1BRESP			(SAXIGP0BRESP	),
	.SAXIGP1BVALID			(SAXIGP0BVALID	),
	.SAXIGP1RDATA			(SAXIGP0RDATA	),
	.SAXIGP1RID			(SAXIGP0RID	),
	.SAXIGP1RLAST			(SAXIGP0RLAST	),
	.SAXIGP1RRESP			(SAXIGP0RRESP	),
	.SAXIGP1RVALID			(SAXIGP0RVALID	),
	.SAXIGP1WREADY			(SAXIGP0WREADY	),
	.SAXIGP0ARESETN			(),
	.SAXIGP0ARREADY			(),
	.SAXIGP0AWREADY			(),
	.SAXIGP0BID			(),
	.SAXIGP0BRESP			(),
	.SAXIGP0BVALID			(),
	.SAXIGP0RDATA			(),
	.SAXIGP0RID			(),
	.SAXIGP0RLAST			(),
	.SAXIGP0RRESP			(),
	.SAXIGP0RVALID			(),
	.SAXIGP0WREADY			(),
	.SAXIHP0ARESETN			(),
	.SAXIHP0ARREADY			(),
	.SAXIHP0AWREADY			(),
	.SAXIHP0BID			(),
	.SAXIHP0BRESP			(),
	.SAXIHP0BVALID			(),
	.SAXIHP0RACOUNT			(),
	.SAXIHP0RCOUNT			(),
	.SAXIHP0RDATA			(),
	.SAXIHP0RID			(),
	.SAXIHP0RLAST			(),
	.SAXIHP0RRESP			(),
	.SAXIHP0RVALID			(),
	.SAXIHP0WACOUNT			(),
	.SAXIHP0WCOUNT			(),
	.SAXIHP0WREADY			(),
	.SAXIHP1ARESETN			(),
	.SAXIHP1ARREADY			(),
	.SAXIHP1AWREADY			(),
	.SAXIHP1BID			(),
	.SAXIHP1BRESP			(),
	.SAXIHP1BVALID			(),
	.SAXIHP1RACOUNT			(),
	.SAXIHP1RCOUNT			(),
	.SAXIHP1RDATA			(),
	.SAXIHP1RID			(),
	.SAXIHP1RLAST			(),
	.SAXIHP1RRESP			(),
	.SAXIHP1RVALID			(),
	.SAXIHP1WACOUNT			(),
	.SAXIHP1WCOUNT			(),
	.SAXIHP1WREADY			(),
	.SAXIHP2ARESETN			(),
	.SAXIHP2ARREADY			(),
	.SAXIHP2AWREADY			(),
	.SAXIHP2BID			(),
	.SAXIHP2BRESP			(),
	.SAXIHP2BVALID			(),
	.SAXIHP2RACOUNT			(),
	.SAXIHP2RCOUNT			(),
	.SAXIHP2RDATA			(),
	.SAXIHP2RID			(),
	.SAXIHP2RLAST			(),
	.SAXIHP2RRESP			(),
	.SAXIHP2RVALID			(),
	.SAXIHP2WACOUNT			(),
	.SAXIHP2WCOUNT			(),
	.SAXIHP2WREADY			(),
	.SAXIHP3ARESETN			(),
	.SAXIHP3ARREADY			(),
	.SAXIHP3AWREADY			(),
	.SAXIHP3BID			(),
	.SAXIHP3BRESP			(),
	.SAXIHP3BVALID			(),
	.SAXIHP3RACOUNT			(),
	.SAXIHP3RCOUNT			(),
	.SAXIHP3RDATA			(),
	.SAXIHP3RID			(),
	.SAXIHP3RLAST			(),
	.SAXIHP3RRESP			(),
	.SAXIHP3RVALID			(),
	.SAXIHP3WACOUNT			(),
	.SAXIHP3WCOUNT			(),
	.SAXIHP3WREADY			(),
	.DDRA				(),
	.DDRBA				(),
	.DDRCASB			(),
	.DDRCKE				(),
	.DDRCKN				(),
	.DDRCKP				(),
	.DDRCSB				(),
	.DDRDM				(),
	.DDRDQ				(),
	.DDRDQSN			(),
	.DDRDQSP			(),
	.DDRDRSTB			(),
	.DDRODT				(),
	.DDRRASB			(),
	.DDRVRN				(),
	.DDRVRP				(),
	.DDRWEB				(),
	.MIO				(),
	.PSCLK				(),
	.PSPORB				(),
	.PSSRSTB			(),
	.DDRARB				(),
	.DMA0ACLK			(),
	.DMA0DAREADY			(),
	.DMA0DRLAST			(),
	.DMA0DRTYPE			(),
	.DMA0DRVALID			(),
	.DMA1ACLK			(),
	.DMA1DAREADY			(),
	.DMA1DRLAST			(),
	.DMA1DRTYPE			(),
	.DMA1DRVALID			(),
	.DMA2ACLK			(),
	.DMA2DAREADY			(),
	.DMA2DRLAST			(),
	.DMA2DRTYPE			(),
	.DMA2DRVALID			(),
	.DMA3ACLK			(),
	.DMA3DAREADY			(),
	.DMA3DRLAST			(),
	.DMA3DRTYPE			(),
	.DMA3DRVALID			(),
	.EMIOCAN0PHYRX			(),
	.EMIOCAN1PHYRX			(),
	.EMIOENET0EXTINTIN		(),
	.EMIOENET0GMIICOL		(),
	.EMIOENET0GMIICRS		(),
	.EMIOENET0GMIIRXCLK		(),
	.EMIOENET0GMIIRXD		(),
	.EMIOENET0GMIIRXDV		(),
	.EMIOENET0GMIIRXER		(),
	.EMIOENET0GMIITXCLK		(),
	.EMIOENET0MDIOI			(),
	.EMIOENET1EXTINTIN		(),
	.EMIOENET1GMIICOL		(),
	.EMIOENET1GMIICRS		(),
	.EMIOENET1GMIIRXCLK		(),
	.EMIOENET1GMIIRXD		(),
	.EMIOENET1GMIIRXDV		(),
	.EMIOENET1GMIIRXER		(),
	.EMIOENET1GMIITXCLK		(),
	.EMIOENET1MDIOI			(),
	.EMIOGPIOI			(),
	.EMIOI2C0SCLI			(),
	.EMIOI2C0SDAI			(),
	.EMIOI2C1SCLI			(),
	.EMIOI2C1SDAI			(),
	.EMIOPJTAGTCK			(),
	.EMIOPJTAGTDI			(),
	.EMIOPJTAGTMS			(),
	.EMIOSDIO0CDN			(),
	.EMIOSDIO0CLKFB			(),
	.EMIOSDIO0CMDI			(),
	.EMIOSDIO0DATAI			(),
	.EMIOSDIO0WP			(),
	.EMIOSDIO1CDN			(),
	.EMIOSDIO1CLKFB			(),
	.EMIOSDIO1CMDI			(),
	.EMIOSDIO1DATAI			(),
	.EMIOSDIO1WP			(),
	.EMIOSPI0MI			(),
	.EMIOSPI0SCLKI			(),
	.EMIOSPI0SI			(),
	.EMIOSPI0SSIN			(),
	.EMIOSPI1MI			(),
	.EMIOSPI1SCLKI			(),
	.EMIOSPI1SI			(),
	.EMIOSPI1SSIN			(),
	.EMIOSRAMINTIN			(),
	.EMIOTRACECLK			(),
	.EMIOTTC0CLKI			(),
	.EMIOTTC1CLKI			(),
	.EMIOUART0CTSN			(),
	.EMIOUART0DCDN			(),
	.EMIOUART0DSRN			(),
	.EMIOUART0RIN			(),
	.EMIOUART0RX			(),
	.EMIOUART1CTSN			(),
	.EMIOUART1DCDN			(),
	.EMIOUART1DSRN			(),
	.EMIOUART1RIN			(),
	.EMIOUART1RX			(),
	.EMIOUSB0VBUSPWRFAULT		(1'b0),
	.EMIOUSB1VBUSPWRFAULT		(1'b0),
	.EMIOWDTCLKI			(),
	.EVENTEVENTI			(),
	.FCLKCLKTRIGN			(),
	.FPGAIDLEN			(),
	.FTMDTRACEINATID		(),
	.FTMDTRACEINCLOCK		(),
	.FTMDTRACEINDATA		(),
	.FTMDTRACEINVALID		(),
	.FTMTF2PDEBUG			(),
	.FTMTF2PTRIG			(),
	.FTMTP2FTRIGACK			(),
	.IRQF2P				(irqf2p),
	.MAXIGP0ACLK			(MAXIGP0ACLK),
	.MAXIGP0ARREADY			(MAXIGP0ARREADY	),
	.MAXIGP0AWREADY			(MAXIGP0AWREADY	),
	.MAXIGP0BID			(MAXIGP0BID),
	.MAXIGP0BRESP			(MAXIGP0BRESP	),
	.MAXIGP0BVALID			(MAXIGP0BVALID	),
	.MAXIGP0RDATA			(MAXIGP0RDATA	),
	.MAXIGP0RID			(MAXIGP0RID),
	.MAXIGP0RLAST			(1'b1),
	.MAXIGP0RRESP			(MAXIGP0RRESP	),
	.MAXIGP0RVALID			(MAXIGP0RVALID	),
	.MAXIGP0WREADY			(MAXIGP0WREADY	),
	.MAXIGP1ACLK			(),
	.MAXIGP1ARREADY			(),
	.MAXIGP1AWREADY			(),
	.MAXIGP1BID			(),
	.MAXIGP1BRESP			(),
	.MAXIGP1BVALID			(),
	.MAXIGP1RDATA			(),
	.MAXIGP1RID			(),
	.MAXIGP1RLAST			(),
	.MAXIGP1RRESP			(),
	.MAXIGP1RVALID			(),
	.MAXIGP1WREADY			(),
	.SAXIACPACLK			(),
	.SAXIACPARADDR			(),
	.SAXIACPARBURST			(),
	.SAXIACPARCACHE			(),
	.SAXIACPARID			(),
	.SAXIACPARLEN			(),
	.SAXIACPARLOCK			(),
	.SAXIACPARPROT			(),
	.SAXIACPARQOS			(),
	.SAXIACPARSIZE			(),
	.SAXIACPARUSER			(),
	.SAXIACPARVALID			(),
	.SAXIACPAWADDR			(),
	.SAXIACPAWBURST			(),
	.SAXIACPAWCACHE			(),
	.SAXIACPAWID			(),
	.SAXIACPAWLEN			(),
	.SAXIACPAWLOCK			(),
	.SAXIACPAWPROT			(),
	.SAXIACPAWQOS			(),
	.SAXIACPAWSIZE			(),
	.SAXIACPAWUSER			(),
	.SAXIACPAWVALID			(),
	.SAXIACPBREADY			(),
	.SAXIACPRREADY			(),
	.SAXIACPWDATA			(),
	.SAXIACPWID			(),
	.SAXIACPWLAST			(),
	.SAXIACPWSTRB			(),
	.SAXIACPWVALID			(),
	/* SAXI GP0 inputs */
	.SAXIGP1ACLK			(SAXIGP0ACLK	),
	.SAXIGP1ARADDR			(SAXIGP0ARADDR	),
	.SAXIGP1ARBURST			(SAXIGP0ARBURST	),
	.SAXIGP1ARCACHE			(SAXIGP0ARCACHE	),
	.SAXIGP1ARID			(SAXIGP0ARID	),
	.SAXIGP1ARLEN			(SAXIGP0ARLEN	),
	.SAXIGP1ARLOCK			(SAXIGP0ARLOCK	),
	.SAXIGP1ARPROT			(SAXIGP0ARPROT	),
	.SAXIGP1ARQOS			(SAXIGP0ARQOS	),
	.SAXIGP1ARSIZE			(SAXIGP0ARSIZE	),
	.SAXIGP1ARVALID			(SAXIGP0ARVALID	),
	.SAXIGP1AWADDR			(SAXIGP0AWADDR	),
	.SAXIGP1AWBURST			(SAXIGP0AWBURST	),
	.SAXIGP1AWCACHE			(SAXIGP0AWCACHE	),
	.SAXIGP1AWID			(SAXIGP0AWID	),
	.SAXIGP1AWLEN			(SAXIGP0AWLEN	),
	.SAXIGP1AWLOCK			(SAXIGP0AWLOCK	),
	.SAXIGP1AWPROT			(SAXIGP0AWPROT	),
	.SAXIGP1AWQOS			(SAXIGP0AWQOS	),
	.SAXIGP1AWSIZE			(SAXIGP0AWSIZE	),
	.SAXIGP1AWVALID			(SAXIGP0AWVALID	),
	.SAXIGP1BREADY			(SAXIGP0BREADY	),
	.SAXIGP1RREADY			(SAXIGP0RREADY	),
	.SAXIGP1WDATA			(SAXIGP0WDATA	),
	.SAXIGP1WID			(SAXIGP0WID	),
	.SAXIGP1WLAST			(SAXIGP0WLAST	),
	.SAXIGP1WSTRB			(SAXIGP0WSTRB	),
	.SAXIGP1WVALID			(SAXIGP0WVALID	),
	.SAXIGP0ACLK			(),
	.SAXIGP0ARADDR			(),
	.SAXIGP0ARBURST			(),
	.SAXIGP0ARCACHE			(),
	.SAXIGP0ARID			(),
	.SAXIGP0ARLEN			(),
	.SAXIGP0ARLOCK			(),
	.SAXIGP0ARPROT			(),
	.SAXIGP0ARQOS			(),
	.SAXIGP0ARSIZE			(),
	.SAXIGP0ARVALID			(),
	.SAXIGP0AWADDR			(),
	.SAXIGP0AWBURST			(),
	.SAXIGP0AWCACHE			(),
	.SAXIGP0AWID			(),
	.SAXIGP0AWLEN			(),
	.SAXIGP0AWLOCK			(),
	.SAXIGP0AWPROT			(),
	.SAXIGP0AWQOS			(),
	.SAXIGP0AWSIZE			(),
	.SAXIGP0AWVALID			(),
	.SAXIGP0BREADY			(),
	.SAXIGP0RREADY			(),
	.SAXIGP0WDATA			(),
	.SAXIGP0WID			(),
	.SAXIGP0WLAST			(),
	.SAXIGP0WSTRB			(),
	.SAXIGP0WVALID			(),
	.SAXIHP0ACLK			(),
	.SAXIHP0ARADDR			(),
	.SAXIHP0ARBURST			(),
	.SAXIHP0ARCACHE			(),
	.SAXIHP0ARID			(),
	.SAXIHP0ARLEN			(),
	.SAXIHP0ARLOCK			(),
	.SAXIHP0ARPROT			(),
	.SAXIHP0ARQOS			(),
	.SAXIHP0ARSIZE			(),
	.SAXIHP0ARVALID			(),
	.SAXIHP0AWADDR			(),
	.SAXIHP0AWBURST			(),
	.SAXIHP0AWCACHE			(),
	.SAXIHP0AWID			(),
	.SAXIHP0AWLEN			(),
	.SAXIHP0AWLOCK			(),
	.SAXIHP0AWPROT			(),
	.SAXIHP0AWQOS			(),
	.SAXIHP0AWSIZE			(),
	.SAXIHP0AWVALID			(),
	.SAXIHP0BREADY			(),
	.SAXIHP0RDISSUECAP1EN		(),
	.SAXIHP0RREADY			(),
	.SAXIHP0WDATA			(),
	.SAXIHP0WID			(),
	.SAXIHP0WLAST			(),
	.SAXIHP0WRISSUECAP1EN		(),
	.SAXIHP0WSTRB			(),
	.SAXIHP0WVALID			(),
	.SAXIHP1ACLK			(),
	.SAXIHP1ARADDR			(),
	.SAXIHP1ARBURST			(),
	.SAXIHP1ARCACHE			(),
	.SAXIHP1ARID			(),
	.SAXIHP1ARLEN			(),
	.SAXIHP1ARLOCK			(),
	.SAXIHP1ARPROT			(),
	.SAXIHP1ARQOS			(),
	.SAXIHP1ARSIZE			(),
	.SAXIHP1ARVALID			(),
	.SAXIHP1AWADDR			(),
	.SAXIHP1AWBURST			(),
	.SAXIHP1AWCACHE			(),
	.SAXIHP1AWID			(),
	.SAXIHP1AWLEN			(),
	.SAXIHP1AWLOCK			(),
	.SAXIHP1AWPROT			(),
	.SAXIHP1AWQOS			(),
	.SAXIHP1AWSIZE			(),
	.SAXIHP1AWVALID			(),
	.SAXIHP1BREADY			(),
	.SAXIHP1RDISSUECAP1EN		(),
	.SAXIHP1RREADY			(),
	.SAXIHP1WDATA			(),
	.SAXIHP1WID			(),
	.SAXIHP1WLAST			(),
	.SAXIHP1WRISSUECAP1EN		(),
	.SAXIHP1WSTRB			(),
	.SAXIHP1WVALID			(),
	.SAXIHP2ACLK			(),
	.SAXIHP2ARADDR			(),
	.SAXIHP2ARBURST			(),
	.SAXIHP2ARCACHE			(),
	.SAXIHP2ARID			(),
	.SAXIHP2ARLEN			(),
	.SAXIHP2ARLOCK			(),
	.SAXIHP2ARPROT			(),
	.SAXIHP2ARQOS			(),
	.SAXIHP2ARSIZE			(),
	.SAXIHP2ARVALID			(),
	.SAXIHP2AWADDR			(),
	.SAXIHP2AWBURST			(),
	.SAXIHP2AWCACHE			(),
	.SAXIHP2AWID			(),
	.SAXIHP2AWLEN			(),
	.SAXIHP2AWLOCK			(),
	.SAXIHP2AWPROT			(),
	.SAXIHP2AWQOS			(),
	.SAXIHP2AWSIZE			(),
	.SAXIHP2AWVALID			(),
	.SAXIHP2BREADY			(),
	.SAXIHP2RDISSUECAP1EN		(),
	.SAXIHP2RREADY			(),
	.SAXIHP2WDATA			(),
	.SAXIHP2WID			(),
	.SAXIHP2WLAST			(),
	.SAXIHP2WRISSUECAP1EN		(),
	.SAXIHP2WSTRB			(),
	.SAXIHP2WVALID			(),
	.SAXIHP3ACLK			(),
	.SAXIHP3ARADDR			(),
	.SAXIHP3ARBURST			(),
	.SAXIHP3ARCACHE			(),
	.SAXIHP3ARID			(),
	.SAXIHP3ARLEN			(),
	.SAXIHP3ARLOCK			(),
	.SAXIHP3ARPROT			(),
	.SAXIHP3ARQOS			(),
	.SAXIHP3ARSIZE			(),
	.SAXIHP3ARVALID			(),
	.SAXIHP3AWADDR			(),
	.SAXIHP3AWBURST			(),
	.SAXIHP3AWCACHE			(),
	.SAXIHP3AWID			(),
	.SAXIHP3AWLEN			(),
	.SAXIHP3AWLOCK			(),
	.SAXIHP3AWPROT			(),
	.SAXIHP3AWQOS			(),
	.SAXIHP3AWSIZE			(),
	.SAXIHP3AWVALID			(),
	.SAXIHP3BREADY			(),
	.SAXIHP3RDISSUECAP1EN		(),
	.SAXIHP3RREADY			(),
	.SAXIHP3WDATA			(),
	.SAXIHP3WID			(),
	.SAXIHP3WLAST			(),
	.SAXIHP3WRISSUECAP1EN		(),
	.SAXIHP3WSTRB			(),
	.SAXIHP3WVALID			()
	);

AxiPeriph testSlave (
	.clock(fclk0_bg),
	.reset(reset),
	.io_axi_s0_aw_awaddr(MAXIGP0AWADDR),
	.io_axi_s0_aw_awprot(MAXIGP0AWPROT),
	.io_axi_s0_aw_awvalid(MAXIGP0AWVALID),
	.io_axi_s0_aw_awready(MAXIGP0AWREADY),
	.io_axi_s0_aw_awid(MAXIGP0AWID),
	.io_axi_s0_w_wdata(MAXIGP0WDATA),
	.io_axi_s0_w_wstrb(MAXIGP0WSTRB),
	.io_axi_s0_w_wvalid(MAXIGP0WVALID),
	.io_axi_s0_w_wready(MAXIGP0WREADY),
	.io_axi_s0_w_wid(MAXIGP0WID),
	.io_axi_s0_b_bresp(MAXIGP0BRESP),
	.io_axi_s0_b_bvalid(MAXIGP0BVALID),
	.io_axi_s0_b_bready(MAXIGP0BREADY),
	.io_axi_s0_b_bid(MAXIGP0BID),
	.io_axi_s0_ar_araddr(MAXIGP0ARADDR),
	.io_axi_s0_ar_arprot(MAXIGP0ARPROT),
	.io_axi_s0_ar_arready(MAXIGP0ARREADY),
	.io_axi_s0_ar_arvalid(MAXIGP0ARVALID),
	.io_axi_s0_ar_arid(MAXIGP0ARID),
	.io_axi_s0_r_rdata(MAXIGP0RDATA),
	.io_axi_s0_r_rresp(MAXIGP0RRESP),
	.io_axi_s0_r_rvalid(MAXIGP0RVALID),
	.io_axi_s0_r_rready(MAXIGP0RREADY),
	.io_axi_s0_r_rid(MAXIGP0RID),
	.io_leds(gpios),
	.io_irqOut(testirq_f2p),
	.io_raddr(SAXIGP0ARADDR),
	.io_waddr(SAXIGP0AWADDR),
	.io_rdata(SAXIGP0RDATA),
	.io_wdata(SAXIGP0WDATA)
);

litex_top LitexTop(
	.serial_tx		(tx		),
	.serial_rx		(rx		),
	.cpu_reset		(litex_reset	),
	.clk			(clk125_bg	),
	.clk_out		(fclk0_bg	),
	.s_axi_axi_awready	(SAXIGP0AWREADY	),
	.s_axi_axi_awid		(SAXIGP0AWID	),
	.s_axi_axi_awaddr	(SAXIGP0AWADDR	),
	.s_axi_axi_awlen	(SAXIGP0AWLEN	),
	.s_axi_axi_awsize	(SAXIGP0AWSIZE	),
	.s_axi_axi_awburst	(SAXIGP0AWBURST	),
	.s_axi_axi_awlock	(SAXIGP0AWLOCK	),
	.s_axi_axi_awcache	(SAXIGP0AWCACHE	),
	.s_axi_axi_awprot	(SAXIGP0AWPROT	),
	.s_axi_axi_awqos	(SAXIGP0AWQOS	),
	.s_axi_axi_awvalid	(SAXIGP0AWVALID	),
	.s_axi_axi_wready	(SAXIGP0WREADY	),
	.s_axi_axi_wdata	(SAXIGP0WDATA	),
	.s_axi_axi_wstrb	(SAXIGP0WSTRB	),
	.s_axi_axi_wlast	(SAXIGP0WLAST	),
	.s_axi_axi_wvalid	(SAXIGP0WVALID	),
	.s_axi_axi_bid		(SAXIGP0BID	),
	.s_axi_axi_bresp	(SAXIGP0BRESP	),
	.s_axi_axi_bvalid	(SAXIGP0BVALID	),
	.s_axi_axi_bready	(SAXIGP0BREADY	),
	.s_axi_axi_arready	(SAXIGP0ARREADY	),
	.s_axi_axi_arid		(SAXIGP0ARID	),
	.s_axi_axi_araddr	(SAXIGP0ARADDR	),
	.s_axi_axi_arlen	(SAXIGP0ARLEN	),
	.s_axi_axi_arsize	(SAXIGP0ARSIZE	),
	.s_axi_axi_arburst	(SAXIGP0ARBURST	),
	.s_axi_axi_arlock	(SAXIGP0ARLOCK	),
	.s_axi_axi_arcache	(SAXIGP0ARCACHE	),
	.s_axi_axi_arprot	(SAXIGP0ARPROT	),
	.s_axi_axi_arqos	(SAXIGP0ARQOS	),
	.s_axi_axi_arvalid	(SAXIGP0ARVALID	),
	.s_axi_axi_rresp	(SAXIGP0RRESP	),
	.s_axi_axi_rvalid	(SAXIGP0RVALID	),
	.s_axi_axi_rdata	(SAXIGP0RDATA	),
	.s_axi_axi_rlast	(SAXIGP0RLAST	),
	.s_axi_axi_rid		(SAXIGP0RID	),
	.s_axi_axi_rready	(SAXIGP0RREADY	)
);
endmodule
