module alert_handler (
	clk_i,
	rst_ni,
	tl_i,
	tl_o,
	intr_classa_o,
	intr_classb_o,
	intr_classc_o,
	intr_classd_o,
	crashdump_o,
	entropy_i,
	alert_tx_i,
	alert_rx_o,
	esc_rx_i,
	esc_tx_o
);
	parameter signed [31:0] alert_handler_reg_pkg_AccuCntDw = 16;
	parameter [alert_handler_reg_pkg_NAlerts - 1:0] alert_handler_reg_pkg_AsyncOn = 1'b0;
	parameter signed [31:0] alert_handler_reg_pkg_CLASS_DW = 2;
	parameter signed [31:0] alert_handler_reg_pkg_EscCntDw = 32;
	parameter signed [31:0] alert_handler_reg_pkg_LfsrSeed = 2147483647;
	parameter signed [31:0] alert_handler_reg_pkg_NAlerts = 1;
	parameter signed [31:0] alert_handler_reg_pkg_N_CLASSES = 4;
	parameter signed [31:0] alert_handler_reg_pkg_N_ESC_SEV = 4;
	parameter signed [31:0] alert_handler_reg_pkg_N_LOC_ALERT = 4;
	parameter signed [31:0] alert_handler_reg_pkg_N_PHASES = 4;
	parameter signed [31:0] alert_handler_reg_pkg_PHASE_DW = 2;
	parameter signed [31:0] alert_handler_reg_pkg_PING_CNT_DW = 24;
	localparam top_pkg_TL_AIW = 8;
	localparam top_pkg_TL_AW = 32;
	localparam top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam top_pkg_TL_DIW = 1;
	localparam top_pkg_TL_DUW = 16;
	localparam top_pkg_TL_DW = 32;
	localparam top_pkg_TL_SZW = $clog2($clog2(32 >> 3) + 1);
	localparam [31:0] NAlerts = alert_handler_reg_pkg_NAlerts;
	localparam [31:0] EscCntDw = alert_handler_reg_pkg_EscCntDw;
	localparam [31:0] AccuCntDw = alert_handler_reg_pkg_AccuCntDw;
	localparam [31:0] LfsrSeed = alert_handler_reg_pkg_LfsrSeed;
	localparam [NAlerts - 1:0] AsyncOn = alert_handler_reg_pkg_AsyncOn;
	localparam [31:0] N_CLASSES = alert_handler_reg_pkg_N_CLASSES;
	localparam [31:0] N_ESC_SEV = alert_handler_reg_pkg_N_ESC_SEV;
	localparam [31:0] N_PHASES = alert_handler_reg_pkg_N_PHASES;
	localparam [31:0] N_LOC_ALERT = alert_handler_reg_pkg_N_LOC_ALERT;
	localparam [31:0] PING_CNT_DW = alert_handler_reg_pkg_PING_CNT_DW;
	localparam [31:0] PHASE_DW = alert_handler_reg_pkg_PHASE_DW;
	localparam [31:0] CLASS_DW = alert_handler_reg_pkg_CLASS_DW;
	localparam [2:0] Idle = 3'b000;
	localparam [2:0] Timeout = 3'b001;
	localparam [2:0] Terminal = 3'b011;
	localparam [2:0] Phase0 = 3'b100;
	localparam [2:0] Phase1 = 3'b101;
	localparam [2:0] Phase2 = 3'b110;
	localparam [2:0] Phase3 = 3'b111;
	input clk_i;
	input rst_ni;
	input wire [((((((7 + ((top_pkg_TL_SZW - 1) >= 0 ? top_pkg_TL_SZW : 2 - top_pkg_TL_SZW)) + top_pkg_TL_AIW) + top_pkg_TL_AW) + ((top_pkg_TL_DBW - 1) >= 0 ? top_pkg_TL_DBW : 2 - top_pkg_TL_DBW)) + top_pkg_TL_DW) + 17) - 1:0] tl_i;
	output wire [((((((7 + ((top_pkg_TL_SZW - 1) >= 0 ? top_pkg_TL_SZW : 2 - top_pkg_TL_SZW)) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + top_pkg_TL_DUW) + 2) - 1:0] tl_o;
	output wire intr_classa_o;
	output wire intr_classb_o;
	output wire intr_classc_o;
	output wire intr_classd_o;
	output wire [((((((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT)) + (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1)) + (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1)) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1)) - 1:0] crashdump_o;
	input entropy_i;
	input wire [((NAlerts - 1) >= 0 ? (NAlerts * 2) + -1 : ((2 - NAlerts) * 2) + (((NAlerts - 1) * 2) - 1)):((NAlerts - 1) >= 0 ? 0 : (NAlerts - 1) * 2)] alert_tx_i;
	output wire [((NAlerts - 1) >= 0 ? (NAlerts * 4) + -1 : ((2 - NAlerts) * 4) + (((NAlerts - 1) * 4) - 1)):((NAlerts - 1) >= 0 ? 0 : (NAlerts - 1) * 4)] alert_rx_o;
	input wire [((N_ESC_SEV - 1) >= 0 ? (N_ESC_SEV * 2) + -1 : ((2 - N_ESC_SEV) * 2) + (((N_ESC_SEV - 1) * 2) - 1)):((N_ESC_SEV - 1) >= 0 ? 0 : (N_ESC_SEV - 1) * 2)] esc_rx_i;
	output wire [((N_ESC_SEV - 1) >= 0 ? (N_ESC_SEV * 2) + -1 : ((2 - N_ESC_SEV) * 2) + (((N_ESC_SEV - 1) * 2) - 1)):((N_ESC_SEV - 1) >= 0 ? 0 : (N_ESC_SEV - 1) * 2)] esc_tx_o;
	wire [N_CLASSES - 1:0] irq;
	wire [((((((((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT)) + ((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES)) + ((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES)) + (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1)) + (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1)) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1)) - 1:0] hw2reg_wrap;
	wire [((((((((((((1 + ((PING_CNT_DW - 1) >= 0 ? PING_CNT_DW : 2 - PING_CNT_DW)) + ((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT)) + (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1)) + ((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts)) + (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1)) + ((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES)) + ((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES)) + (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1)) + (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1)) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1)) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1)) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)) - 1:0] reg2hw_wrap;
	assign {intr_classd_o, intr_classc_o, intr_classb_o, intr_classa_o} = irq;
	alert_handler_reg_wrap i_reg_wrap(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_i(tl_i),
		.tl_o(tl_o),
		.irq_o(irq),
		.crashdump_o(crashdump_o),
		.hw2reg_wrap(hw2reg_wrap),
		.reg2hw_wrap(reg2hw_wrap)
	);
	wire [N_LOC_ALERT - 1:0] loc_alert_trig;
	wire [NAlerts - 1:0] alert_ping_en;
	wire [NAlerts - 1:0] alert_ping_ok;
	wire [N_ESC_SEV - 1:0] esc_ping_en;
	wire [N_ESC_SEV - 1:0] esc_ping_ok;
	alert_handler_ping_timer i_ping_timer(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.entropy_i(entropy_i),
		.en_i(reg2hw_wrap[1 + (((PING_CNT_DW - 1) >= 0 ? PING_CNT_DW : 2 - PING_CNT_DW) + (((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + ((((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))))))))))]),
		.alert_en_i(reg2hw_wrap[((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))))))-:((((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))))))) >= ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)))))))) ? ((((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))))))) - ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1))))))))) + 1 : (((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)))))))) - (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))))))))) + 1)]),
		.ping_timeout_cyc_i(reg2hw_wrap[((PING_CNT_DW - 1) >= 0 ? PING_CNT_DW : 2 - PING_CNT_DW) + (((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + ((((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))))))))))-:((((PING_CNT_DW - 1) >= 0 ? PING_CNT_DW : 2 - PING_CNT_DW) + (((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + ((((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))))))))))) >= (((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + ((((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1))))))))))) ? ((((PING_CNT_DW - 1) >= 0 ? PING_CNT_DW : 2 - PING_CNT_DW) + (((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + ((((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))))))))))) - (((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + ((((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)))))))))))) + 1 : ((((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + ((((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1))))))))))) - (((PING_CNT_DW - 1) >= 0 ? PING_CNT_DW : 2 - PING_CNT_DW) + (((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + ((((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))))))))))) + 1)]),
		.wait_cyc_mask_i(sv2v_cast_3E03F(24'hFFFFFF)),
		.alert_ping_en_o(alert_ping_en),
		.esc_ping_en_o(esc_ping_en),
		.alert_ping_ok_i(alert_ping_ok),
		.esc_ping_ok_i(esc_ping_ok),
		.alert_ping_fail_o(loc_alert_trig[0]),
		.esc_ping_fail_o(loc_alert_trig[1])
	);
	wire [NAlerts - 1:0] alert_integfail;
	wire [NAlerts - 1:0] alert_trig;
	generate
		genvar k;
		for (k = 0; k < NAlerts; k = k + 1) begin : gen_alerts
			prim_alert_receiver #(.AsyncOn(AsyncOn[k])) i_alert_receiver(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.ping_en_i(alert_ping_en[k]),
				.ping_ok_o(alert_ping_ok[k]),
				.integ_fail_o(alert_integfail[k]),
				.alert_o(alert_trig[k]),
				.alert_rx_o(alert_rx_o[((NAlerts - 1) >= 0 ? k : 0 - (k - (NAlerts - 1))) * 4+:4]),
				.alert_tx_i(alert_tx_i[((NAlerts - 1) >= 0 ? k : 0 - (k - (NAlerts - 1))) * 2+:2])
			);
		end
	endgenerate
	assign loc_alert_trig[2] = |(reg2hw_wrap[((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))))))-:((((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))))))) >= ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)))))))) ? ((((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))))))) - ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1))))))))) + 1 : (((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)))))))) - (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))))))))) + 1)] & alert_integfail);
	alert_handler_class i_class(
		.alert_trig_i(alert_trig),
		.loc_alert_trig_i(loc_alert_trig),
		.alert_en_i(reg2hw_wrap[((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))))))-:((((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))))))) >= ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)))))))) ? ((((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))))))) - ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1))))))))) + 1 : (((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)))))))) - (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))))))))) + 1)]),
		.loc_alert_en_i(reg2hw_wrap[((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + ((((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))))))))-:((((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + ((((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))))))))) >= ((((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)))))))))) ? ((((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + ((((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))))))))) - ((((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1))))))))))) + 1 : (((((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)))))))))) - (((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + ((((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))))))))))) + 1)]),
		.alert_class_i(reg2hw_wrap[(((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))))))-:(((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))))))) >= (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1))))))) ? (((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))))))) - (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)))))))) + 1 : ((((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1))))))) - ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))))))) + 1)]),
		.loc_alert_class_i(reg2hw_wrap[(((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))))))))-:(((((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))))))))) >= (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1))))))))) ? (((((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))))))))) - (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)))))))))) + 1 : ((((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1))))))))) - ((((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))))))))) + 1)]),
		.alert_cause_o(hw2reg_wrap[((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + (((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))))))-:((((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + (((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))))))) >= (((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1)))))) ? ((((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + (((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))))))) - (((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1))))))) + 1 : ((((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1)))))) - (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + (((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1)))))))) + 1)]),
		.loc_alert_cause_o(hw2reg_wrap[((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1)))))-:((((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1)))))) >= (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1))))) ? ((((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1)))))) - (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1)))))) + 1 : ((((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1))))) - (((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))))))) + 1)]),
		.class_trig_o(hw2reg_wrap[((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))))-:((((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))))) >= (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1)))) ? ((((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))))) - (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1))))) + 1 : ((((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1)))) - (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1)))))) + 1)])
	);
	wire [N_CLASSES - 1:0] class_accum_trig;
	wire [((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))):((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))] class_esc_sig_en;
	generate
		for (k = 0; k < N_CLASSES; k = k + 1) begin : gen_classes
			alert_handler_accu i_accu(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.class_en_i(reg2hw_wrap[((N_CLASSES - 1) >= 0 ? (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))))) - ((N_CLASSES - 1) - k) : (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)))))) + (0 - k))]),
				.clr_i(reg2hw_wrap[((N_CLASSES - 1) >= 0 ? (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))))) - ((N_CLASSES - 1) - k) : ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1))))) + (0 - k))]),
				.class_trig_i(hw2reg_wrap[((N_CLASSES - 1) >= 0 ? (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))))) - ((N_CLASSES - 1) - k) : (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1)))) + (0 - k))]),
				.thresh_i(reg2hw_wrap[(((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))) - (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - (((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) + (((N_CLASSES - 1) >= 0 ? k : 0 - (k - (N_CLASSES - 1))) * ((AccuCntDw - 1) >= 0 ? AccuCntDw : 2 - AccuCntDw)))) : ((((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)))) + (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - (((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) + (((N_CLASSES - 1) >= 0 ? k : 0 - (k - (N_CLASSES - 1))) * ((AccuCntDw - 1) >= 0 ? AccuCntDw : 2 - AccuCntDw))))) - ((AccuCntDw - 1) >= 0 ? AccuCntDw : 2 - AccuCntDw)) + 1)+:((AccuCntDw - 1) >= 0 ? AccuCntDw : 2 - AccuCntDw)]),
				.accu_cnt_o(hw2reg_wrap[(((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))) - (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - (((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) + (((N_CLASSES - 1) >= 0 ? k : 0 - (k - (N_CLASSES - 1))) * ((AccuCntDw - 1) >= 0 ? AccuCntDw : 2 - AccuCntDw)))) : ((((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1)) + (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - (((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) + (((N_CLASSES - 1) >= 0 ? k : 0 - (k - (N_CLASSES - 1))) * ((AccuCntDw - 1) >= 0 ? AccuCntDw : 2 - AccuCntDw))))) - ((AccuCntDw - 1) >= 0 ? AccuCntDw : 2 - AccuCntDw)) + 1)+:((AccuCntDw - 1) >= 0 ? AccuCntDw : 2 - AccuCntDw)]),
				.accu_trig_o(class_accum_trig[k])
			);
			alert_handler_esc_timer i_esc_timer(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.en_i(reg2hw_wrap[((N_CLASSES - 1) >= 0 ? (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))))) - ((N_CLASSES - 1) - k) : (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)))))) + (0 - k))]),
				.clr_i(reg2hw_wrap[((N_CLASSES - 1) >= 0 ? (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))))) - ((N_CLASSES - 1) - k) : ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1))))) + (0 - k))]),
				.timeout_en_i(irq[k]),
				.accum_trig_i(class_accum_trig[k]),
				.timeout_cyc_i(reg2hw_wrap[(((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))) - (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - (((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? k : 0 - (k - (N_CLASSES - 1))) * ((EscCntDw - 1) >= 0 ? EscCntDw : 2 - EscCntDw)))) : (((((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1))) + (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - (((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? k : 0 - (k - (N_CLASSES - 1))) * ((EscCntDw - 1) >= 0 ? EscCntDw : 2 - EscCntDw))))) - ((EscCntDw - 1) >= 0 ? EscCntDw : 2 - EscCntDw)) + 1)+:((EscCntDw - 1) >= 0 ? EscCntDw : 2 - EscCntDw)]),
				.esc_en_i(reg2hw_wrap[(((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - (((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) + (((N_CLASSES - 1) >= 0 ? k : 0 - (k - (N_CLASSES - 1))) * ((N_ESC_SEV - 1) >= 0 ? N_ESC_SEV : 2 - N_ESC_SEV)))) : ((((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - (((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) + (((N_CLASSES - 1) >= 0 ? k : 0 - (k - (N_CLASSES - 1))) * ((N_ESC_SEV - 1) >= 0 ? N_ESC_SEV : 2 - N_ESC_SEV))))) - ((N_ESC_SEV - 1) >= 0 ? N_ESC_SEV : 2 - N_ESC_SEV)) + 1)+:((N_ESC_SEV - 1) >= 0 ? N_ESC_SEV : 2 - N_ESC_SEV)]),
				.esc_map_i(reg2hw_wrap[((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1) - ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((PHASE_DW - 1) >= 0 ? 0 : PHASE_DW - 1) + (((PHASE_DW - 1) >= 0 ? PHASE_DW : 2 - PHASE_DW) * (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) + (((N_CLASSES - 1) >= 0 ? k : 0 - (k - (N_CLASSES - 1))) * ((N_ESC_SEV - 1) >= 0 ? N_ESC_SEV : 2 - N_ESC_SEV)) : (((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) + (((N_CLASSES - 1) >= 0 ? k : 0 - (k - (N_CLASSES - 1))) * ((N_ESC_SEV - 1) >= 0 ? N_ESC_SEV : 2 - N_ESC_SEV))) + (((N_ESC_SEV - 1) >= 0 ? N_ESC_SEV : 2 - N_ESC_SEV) - 1)) : ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) + (((N_CLASSES - 1) >= 0 ? k : 0 - (k - (N_CLASSES - 1))) * ((N_ESC_SEV - 1) >= 0 ? N_ESC_SEV : 2 - N_ESC_SEV)) : (((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) + (((N_CLASSES - 1) >= 0 ? k : 0 - (k - (N_CLASSES - 1))) * ((N_ESC_SEV - 1) >= 0 ? N_ESC_SEV : 2 - N_ESC_SEV))) + (((N_ESC_SEV - 1) >= 0 ? N_ESC_SEV : 2 - N_ESC_SEV) - 1)) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))))))) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((PHASE_DW - 1) >= 0 ? 0 : PHASE_DW - 1) + (((PHASE_DW - 1) >= 0 ? PHASE_DW : 2 - PHASE_DW) * (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) + (((N_CLASSES - 1) >= 0 ? k : 0 - (k - (N_CLASSES - 1))) * ((N_ESC_SEV - 1) >= 0 ? N_ESC_SEV : 2 - N_ESC_SEV)) : (((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) + (((N_CLASSES - 1) >= 0 ? k : 0 - (k - (N_CLASSES - 1))) * ((N_ESC_SEV - 1) >= 0 ? N_ESC_SEV : 2 - N_ESC_SEV))) + (((N_ESC_SEV - 1) >= 0 ? N_ESC_SEV : 2 - N_ESC_SEV) - 1)) : ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) + (((N_CLASSES - 1) >= 0 ? k : 0 - (k - (N_CLASSES - 1))) * ((N_ESC_SEV - 1) >= 0 ? N_ESC_SEV : 2 - N_ESC_SEV)) : (((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) + (((N_CLASSES - 1) >= 0 ? k : 0 - (k - (N_CLASSES - 1))) * ((N_ESC_SEV - 1) >= 0 ? N_ESC_SEV : 2 - N_ESC_SEV))) + (((N_ESC_SEV - 1) >= 0 ? N_ESC_SEV : 2 - N_ESC_SEV) - 1)) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))))))) - (((PHASE_DW - 1) >= 0 ? PHASE_DW : 2 - PHASE_DW) * ((N_ESC_SEV - 1) >= 0 ? N_ESC_SEV : 2 - N_ESC_SEV))) + 1)+:((PHASE_DW - 1) >= 0 ? PHASE_DW : 2 - PHASE_DW) * ((N_ESC_SEV - 1) >= 0 ? N_ESC_SEV : 2 - N_ESC_SEV)]),
				.phase_cyc_i(reg2hw_wrap[((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))) - ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) + (((EscCntDw - 1) >= 0 ? EscCntDw : 2 - EscCntDw) * (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) + (((N_CLASSES - 1) >= 0 ? k : 0 - (k - (N_CLASSES - 1))) * ((N_PHASES - 1) >= 0 ? N_PHASES : 2 - N_PHASES)) : (((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) + (((N_CLASSES - 1) >= 0 ? k : 0 - (k - (N_CLASSES - 1))) * ((N_PHASES - 1) >= 0 ? N_PHASES : 2 - N_PHASES))) + (((N_PHASES - 1) >= 0 ? N_PHASES : 2 - N_PHASES) - 1)) : ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) + (((N_CLASSES - 1) >= 0 ? k : 0 - (k - (N_CLASSES - 1))) * ((N_PHASES - 1) >= 0 ? N_PHASES : 2 - N_PHASES)) : (((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) + (((N_CLASSES - 1) >= 0 ? k : 0 - (k - (N_CLASSES - 1))) * ((N_PHASES - 1) >= 0 ? N_PHASES : 2 - N_PHASES))) + (((N_PHASES - 1) >= 0 ? N_PHASES : 2 - N_PHASES) - 1)) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))))))) : ((((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) + (((EscCntDw - 1) >= 0 ? EscCntDw : 2 - EscCntDw) * (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) + (((N_CLASSES - 1) >= 0 ? k : 0 - (k - (N_CLASSES - 1))) * ((N_PHASES - 1) >= 0 ? N_PHASES : 2 - N_PHASES)) : (((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) + (((N_CLASSES - 1) >= 0 ? k : 0 - (k - (N_CLASSES - 1))) * ((N_PHASES - 1) >= 0 ? N_PHASES : 2 - N_PHASES))) + (((N_PHASES - 1) >= 0 ? N_PHASES : 2 - N_PHASES) - 1)) : ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) + (((N_CLASSES - 1) >= 0 ? k : 0 - (k - (N_CLASSES - 1))) * ((N_PHASES - 1) >= 0 ? N_PHASES : 2 - N_PHASES)) : (((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) + (((N_CLASSES - 1) >= 0 ? k : 0 - (k - (N_CLASSES - 1))) * ((N_PHASES - 1) >= 0 ? N_PHASES : 2 - N_PHASES))) + (((N_PHASES - 1) >= 0 ? N_PHASES : 2 - N_PHASES) - 1)) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))))))))) - (((EscCntDw - 1) >= 0 ? EscCntDw : 2 - EscCntDw) * ((N_PHASES - 1) >= 0 ? N_PHASES : 2 - N_PHASES))) + 1)+:((EscCntDw - 1) >= 0 ? EscCntDw : 2 - EscCntDw) * ((N_PHASES - 1) >= 0 ? N_PHASES : 2 - N_PHASES)]),
				.esc_trig_o(hw2reg_wrap[((N_CLASSES - 1) >= 0 ? (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1)))) - ((N_CLASSES - 1) - k) : ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1))) + (0 - k))]),
				.esc_cnt_o(hw2reg_wrap[(((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1)) - (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - (((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? k : 0 - (k - (N_CLASSES - 1))) * ((EscCntDw - 1) >= 0 ? EscCntDw : 2 - EscCntDw)))) : (((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - (((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? k : 0 - (k - (N_CLASSES - 1))) * ((EscCntDw - 1) >= 0 ? EscCntDw : 2 - EscCntDw))))) - ((EscCntDw - 1) >= 0 ? EscCntDw : 2 - EscCntDw)) + 1)+:((EscCntDw - 1) >= 0 ? EscCntDw : 2 - EscCntDw)]),
				.esc_state_o(hw2reg_wrap[(((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1) - (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - (((N_CLASSES - 1) >= 0 ? k : 0 - (k - (N_CLASSES - 1))) * 3)) : ((((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - (((N_CLASSES - 1) >= 0 ? k : 0 - (k - (N_CLASSES - 1))) * 3)) - 3) + 1)+:3]),
				.esc_sig_en_o(class_esc_sig_en[((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) + (((N_CLASSES - 1) >= 0 ? k : 0 - (k - (N_CLASSES - 1))) * ((N_ESC_SEV - 1) >= 0 ? N_ESC_SEV : 2 - N_ESC_SEV))+:((N_ESC_SEV - 1) >= 0 ? N_ESC_SEV : 2 - N_ESC_SEV)])
			);
		end
	endgenerate
	wire [N_ESC_SEV - 1:0] esc_sig_en;
	wire [N_ESC_SEV - 1:0] esc_integfail;
	wire [((N_ESC_SEV - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? (N_ESC_SEV * N_CLASSES) + -1 : (N_ESC_SEV * (2 - N_CLASSES)) + ((N_CLASSES - 1) - 1)) : ((N_CLASSES - 1) >= 0 ? ((2 - N_ESC_SEV) * N_CLASSES) + (((N_ESC_SEV - 1) * N_CLASSES) - 1) : ((2 - N_ESC_SEV) * (2 - N_CLASSES)) + (((N_CLASSES - 1) + ((N_ESC_SEV - 1) * (2 - N_CLASSES))) - 1))):((N_ESC_SEV - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? 0 : N_CLASSES - 1) : ((N_CLASSES - 1) >= 0 ? (N_ESC_SEV - 1) * N_CLASSES : (N_CLASSES - 1) + ((N_ESC_SEV - 1) * (2 - N_CLASSES))))] esc_sig_en_trsp;
	generate
		genvar j;
		for (k = 0; k < N_ESC_SEV; k = k + 1) begin : gen_esc_sev
			for (j = 0; j < N_CLASSES; j = j + 1) begin : gen_transp
				assign esc_sig_en_trsp[(((N_ESC_SEV - 1) >= 0 ? k : 0 - (k - (N_ESC_SEV - 1))) * ((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES)) + ((N_CLASSES - 1) >= 0 ? j : 0 - (j - (N_CLASSES - 1)))] = class_esc_sig_en[(((N_CLASSES - 1) >= 0 ? j : 0 - (j - (N_CLASSES - 1))) * ((N_ESC_SEV - 1) >= 0 ? N_ESC_SEV : 2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) >= 0 ? k : 0 - (k - (N_ESC_SEV - 1)))];
			end
			assign esc_sig_en[k] = |esc_sig_en_trsp[((N_CLASSES - 1) >= 0 ? 0 : N_CLASSES - 1) + (((N_ESC_SEV - 1) >= 0 ? k : 0 - (k - (N_ESC_SEV - 1))) * ((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES))+:((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES)];
			prim_esc_sender i_esc_sender(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.ping_en_i(esc_ping_en[k]),
				.ping_ok_o(esc_ping_ok[k]),
				.integ_fail_o(esc_integfail[k]),
				.esc_en_i(esc_sig_en[k]),
				.esc_rx_i(esc_rx_i[((N_ESC_SEV - 1) >= 0 ? k : 0 - (k - (N_ESC_SEV - 1))) * 2+:2]),
				.esc_tx_o(esc_tx_o[((N_ESC_SEV - 1) >= 0 ? k : 0 - (k - (N_ESC_SEV - 1))) * 2+:2])
			);
		end
	endgenerate
	assign loc_alert_trig[3] = |esc_integfail;
	function automatic [alert_handler_reg_pkg_PING_CNT_DW - 1:0] sv2v_cast_3E03F;
		input reg [alert_handler_reg_pkg_PING_CNT_DW - 1:0] inp;
		sv2v_cast_3E03F = inp;
	endfunction
endmodule
