module alert_handler_reg_wrap (
	clk_i,
	rst_ni,
	tl_i,
	tl_o,
	irq_o,
	crashdump_o,
	hw2reg_wrap,
	reg2hw_wrap
);
	parameter signed [31:0] alert_handler_reg_pkg_AccuCntDw = 16;
	parameter [alert_handler_reg_pkg_NAlerts - 1:0] alert_handler_reg_pkg_AsyncOn = 1'b0;
	parameter signed [31:0] alert_handler_reg_pkg_CLASS_DW = 2;
	parameter signed [31:0] alert_handler_reg_pkg_EscCntDw = 32;
	parameter signed [31:0] alert_handler_reg_pkg_LfsrSeed = 2147483647;
	parameter signed [31:0] alert_handler_reg_pkg_NAlerts = 1;
	parameter signed [31:0] alert_handler_reg_pkg_N_CLASSES = 4;
	parameter signed [31:0] alert_handler_reg_pkg_N_ESC_SEV = 4;
	parameter signed [31:0] alert_handler_reg_pkg_N_LOC_ALERT = 4;
	parameter signed [31:0] alert_handler_reg_pkg_N_PHASES = 4;
	parameter signed [31:0] alert_handler_reg_pkg_PHASE_DW = 2;
	parameter signed [31:0] alert_handler_reg_pkg_PING_CNT_DW = 24;
	localparam top_pkg_TL_AIW = 8;
	localparam top_pkg_TL_AW = 32;
	localparam top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam top_pkg_TL_DIW = 1;
	localparam top_pkg_TL_DUW = 16;
	localparam top_pkg_TL_DW = 32;
	localparam top_pkg_TL_SZW = $clog2($clog2(32 >> 3) + 1);
	localparam [31:0] NAlerts = alert_handler_reg_pkg_NAlerts;
	localparam [31:0] EscCntDw = alert_handler_reg_pkg_EscCntDw;
	localparam [31:0] AccuCntDw = alert_handler_reg_pkg_AccuCntDw;
	localparam [31:0] LfsrSeed = alert_handler_reg_pkg_LfsrSeed;
	localparam [NAlerts - 1:0] AsyncOn = alert_handler_reg_pkg_AsyncOn;
	localparam [31:0] N_CLASSES = alert_handler_reg_pkg_N_CLASSES;
	localparam [31:0] N_ESC_SEV = alert_handler_reg_pkg_N_ESC_SEV;
	localparam [31:0] N_PHASES = alert_handler_reg_pkg_N_PHASES;
	localparam [31:0] N_LOC_ALERT = alert_handler_reg_pkg_N_LOC_ALERT;
	localparam [31:0] PING_CNT_DW = alert_handler_reg_pkg_PING_CNT_DW;
	localparam [31:0] PHASE_DW = alert_handler_reg_pkg_PHASE_DW;
	localparam [31:0] CLASS_DW = alert_handler_reg_pkg_CLASS_DW;
	localparam [2:0] Idle = 3'b000;
	localparam [2:0] Timeout = 3'b001;
	localparam [2:0] Terminal = 3'b011;
	localparam [2:0] Phase0 = 3'b100;
	localparam [2:0] Phase1 = 3'b101;
	localparam [2:0] Phase2 = 3'b110;
	localparam [2:0] Phase3 = 3'b111;
	input clk_i;
	input rst_ni;
	input wire [((((((7 + ((top_pkg_TL_SZW - 1) >= 0 ? top_pkg_TL_SZW : 2 - top_pkg_TL_SZW)) + top_pkg_TL_AIW) + top_pkg_TL_AW) + ((top_pkg_TL_DBW - 1) >= 0 ? top_pkg_TL_DBW : 2 - top_pkg_TL_DBW)) + top_pkg_TL_DW) + 17) - 1:0] tl_i;
	output wire [((((((7 + ((top_pkg_TL_SZW - 1) >= 0 ? top_pkg_TL_SZW : 2 - top_pkg_TL_SZW)) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + top_pkg_TL_DUW) + 2) - 1:0] tl_o;
	output wire [N_CLASSES - 1:0] irq_o;
	output wire [((((((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT)) + (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1)) + (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1)) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1)) - 1:0] crashdump_o;
	input wire [((((((((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT)) + ((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES)) + ((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES)) + (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1)) + (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1)) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1)) - 1:0] hw2reg_wrap;
	output wire [((((((((((((1 + ((PING_CNT_DW - 1) >= 0 ? PING_CNT_DW : 2 - PING_CNT_DW)) + ((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT)) + (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1)) + ((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts)) + (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1)) + ((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES)) + ((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES)) + (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1)) + (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1)) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1)) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1)) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)) - 1:0] reg2hw_wrap;
	wire [N_CLASSES - 1:0] class_autolock_en;
	wire [828:0] reg2hw;
	wire [229:0] hw2reg;
	alert_handler_reg_top i_reg(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_i(tl_i),
		.tl_o(tl_o),
		.reg2hw(reg2hw),
		.hw2reg(hw2reg),
		.devmode_i(1'b1)
	);
	prim_intr_hw #(.Width(1)) i_irq_classa(
		.event_intr_i(hw2reg_wrap[((N_CLASSES - 1) >= 0 ? (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))))) - (N_CLASSES - 1) : ((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1))))]),
		.reg2hw_intr_enable_q_i(reg2hw[824]),
		.reg2hw_intr_test_q_i(reg2hw[820]),
		.reg2hw_intr_test_qe_i(reg2hw[819]),
		.reg2hw_intr_state_q_i(reg2hw[828]),
		.hw2reg_intr_state_de_o(hw2reg[228]),
		.hw2reg_intr_state_d_o(hw2reg[229]),
		.intr_o(irq_o[0])
	);
	prim_intr_hw #(.Width(1)) i_irq_classb(
		.event_intr_i(hw2reg_wrap[((N_CLASSES - 1) >= 0 ? (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))))) - ((N_CLASSES - 1) - 1) : (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1)))) + -1)]),
		.reg2hw_intr_enable_q_i(reg2hw[823]),
		.reg2hw_intr_test_q_i(reg2hw[818]),
		.reg2hw_intr_test_qe_i(reg2hw[817]),
		.reg2hw_intr_state_q_i(reg2hw[827]),
		.hw2reg_intr_state_de_o(hw2reg[226]),
		.hw2reg_intr_state_d_o(hw2reg[227]),
		.intr_o(irq_o[1])
	);
	prim_intr_hw #(.Width(1)) i_irq_classc(
		.event_intr_i(hw2reg_wrap[((N_CLASSES - 1) >= 0 ? (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))))) - ((N_CLASSES - 1) - 2) : (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1)))) + -2)]),
		.reg2hw_intr_enable_q_i(reg2hw[822]),
		.reg2hw_intr_test_q_i(reg2hw[816]),
		.reg2hw_intr_test_qe_i(reg2hw[815]),
		.reg2hw_intr_state_q_i(reg2hw[826]),
		.hw2reg_intr_state_de_o(hw2reg[224]),
		.hw2reg_intr_state_d_o(hw2reg[225]),
		.intr_o(irq_o[2])
	);
	prim_intr_hw #(.Width(1)) i_irq_classd(
		.event_intr_i(hw2reg_wrap[((N_CLASSES - 1) >= 0 ? (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))))) - ((N_CLASSES - 1) - 3) : (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1)))) + -3)]),
		.reg2hw_intr_enable_q_i(reg2hw[821]),
		.reg2hw_intr_test_q_i(reg2hw[814]),
		.reg2hw_intr_test_qe_i(reg2hw[813]),
		.reg2hw_intr_state_q_i(reg2hw[825]),
		.hw2reg_intr_state_de_o(hw2reg[222]),
		.hw2reg_intr_state_d_o(hw2reg[223]),
		.intr_o(irq_o[3])
	);
	generate
		genvar k;
		for (k = 0; k < NAlerts; k = k + 1) begin : gen_alert_cause
			assign hw2reg[220 + ((k * 2) + 1)] = 1'b1;
			assign hw2reg[220 + (k * 2)] = reg2hw[784 + k] | hw2reg_wrap[((NAlerts - 1) >= 0 ? (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + (((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))))))) - ((NAlerts - 1) - k) : (((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1)))))) + (0 - k))];
		end
	endgenerate
	generate
		for (k = 0; k < N_LOC_ALERT; k = k + 1) begin : gen_loc_alert_cause
			assign hw2reg[212 + ((k * 2) + 1)] = 1'b1;
			assign hw2reg[212 + (k * 2)] = reg2hw[768 + k] | hw2reg_wrap[((N_LOC_ALERT - 1) >= 0 ? (((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1)))))) - ((N_LOC_ALERT - 1) - k) : (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1))))) + (0 - k))];
		end
	endgenerate
	assign {hw2reg[52], hw2reg[105], hw2reg[158], hw2reg[211]} = 1'sb0;
	assign {hw2reg[51], hw2reg[104], hw2reg[157], hw2reg[210]} = (hw2reg_wrap[((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1)))-:((((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1)))) >= ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1))) ? ((((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1)))) - ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1)))) + 1 : (((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1))) - (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))))) + 1)] & class_autolock_en) & reg2hw_wrap[((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))))-:((((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))))) >= (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)))))) ? ((((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))))) - (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1))))))) + 1 : ((((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)))))) - (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))))))) + 1)];
	assign {hw2reg[50-:16], hw2reg[103-:16], hw2reg[156-:16], hw2reg[209-:16]} = hw2reg_wrap[(((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))-:(((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))) >= ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1)) ? (((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))) - ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1))) + 1 : (((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1)) - ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1)))) + 1)];
	assign {hw2reg[34-:32], hw2reg[87-:32], hw2reg[140-:32], hw2reg[193-:32]} = hw2reg_wrap[(((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1)-:(((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1)) >= (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) ? (((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1)) - (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1)) + 1 : ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) - ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))) + 1)];
	assign {hw2reg[2-:3], hw2reg[55-:3], hw2reg[108-:3], hw2reg[161-:3]} = hw2reg_wrap[(((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1-:(((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1) >= 0 ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) : 1 - ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))];
	assign reg2hw_wrap[1 + (((PING_CNT_DW - 1) >= 0 ? PING_CNT_DW : 2 - PING_CNT_DW) + (((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + ((((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))))))))))] = ~reg2hw[812];
	generate
		for (k = 0; k < NAlerts; k = k + 1) begin : gen_alert_en_class
			assign reg2hw_wrap[((NAlerts - 1) >= 0 ? (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))))))) - ((NAlerts - 1) - k) : ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)))))))) + (0 - k))] = reg2hw[787 + k];
			assign reg2hw_wrap[(((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))))))) - (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - (((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) + (((NAlerts - 1) >= 0 ? k : 0 - (k - (NAlerts - 1))) * ((CLASS_DW - 1) >= 0 ? CLASS_DW : 2 - CLASS_DW)))) : (((((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1))))))) + (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - (((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) + (((NAlerts - 1) >= 0 ? k : 0 - (k - (NAlerts - 1))) * ((CLASS_DW - 1) >= 0 ? CLASS_DW : 2 - CLASS_DW))))) - ((CLASS_DW - 1) >= 0 ? CLASS_DW : 2 - CLASS_DW)) + 1)+:((CLASS_DW - 1) >= 0 ? CLASS_DW : 2 - CLASS_DW)] = reg2hw[785 + ((k * 2) + 1)-:2];
		end
	endgenerate
	generate
		for (k = 0; k < N_LOC_ALERT; k = k + 1) begin : gen_loc_alert_en_class
			assign reg2hw_wrap[((N_LOC_ALERT - 1) >= 0 ? (((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + ((((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))))))))) - ((N_LOC_ALERT - 1) - k) : ((((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)))))))))) + (0 - k))] = reg2hw[780 + k];
			assign reg2hw_wrap[(((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? ((((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))))))))) - (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - (((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) + (((N_LOC_ALERT - 1) >= 0 ? k : 0 - (k - (N_LOC_ALERT - 1))) * ((CLASS_DW - 1) >= 0 ? CLASS_DW : 2 - CLASS_DW)))) : (((((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1))))))))) + (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - (((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) + (((N_LOC_ALERT - 1) >= 0 ? k : 0 - (k - (N_LOC_ALERT - 1))) * ((CLASS_DW - 1) >= 0 ? CLASS_DW : 2 - CLASS_DW))))) - ((CLASS_DW - 1) >= 0 ? CLASS_DW : 2 - CLASS_DW)) + 1)+:((CLASS_DW - 1) >= 0 ? CLASS_DW : 2 - CLASS_DW)] = reg2hw[772 + ((k * 2) + 1)-:2];
		end
	endgenerate
	assign reg2hw_wrap[((PING_CNT_DW - 1) >= 0 ? PING_CNT_DW : 2 - PING_CNT_DW) + (((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + ((((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))))))))))-:((((PING_CNT_DW - 1) >= 0 ? PING_CNT_DW : 2 - PING_CNT_DW) + (((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + ((((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))))))))))) >= (((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + ((((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1))))))))))) ? ((((PING_CNT_DW - 1) >= 0 ? PING_CNT_DW : 2 - PING_CNT_DW) + (((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + ((((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))))))))))) - (((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + ((((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)))))))))))) + 1 : ((((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + ((((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1))))))))))) - (((PING_CNT_DW - 1) >= 0 ? PING_CNT_DW : 2 - PING_CNT_DW) + (((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + ((((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) >= ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) ? (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))))) + 1 : (((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT - 1) * CLASS_DW : (CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW)))) - ((N_LOC_ALERT - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (N_LOC_ALERT * CLASS_DW) + -1 : (N_LOC_ALERT * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - N_LOC_ALERT) * CLASS_DW) + (((N_LOC_ALERT - 1) * CLASS_DW) - 1) : ((2 - N_LOC_ALERT) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((N_LOC_ALERT - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + ((((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) >= ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) ? (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))))) + 1 : (((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? 0 : CLASS_DW - 1) : ((CLASS_DW - 1) >= 0 ? (NAlerts - 1) * CLASS_DW : (CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW)))) - ((NAlerts - 1) >= 0 ? ((CLASS_DW - 1) >= 0 ? (NAlerts * CLASS_DW) + -1 : (NAlerts * (2 - CLASS_DW)) + ((CLASS_DW - 1) - 1)) : ((CLASS_DW - 1) >= 0 ? ((2 - NAlerts) * CLASS_DW) + (((NAlerts - 1) * CLASS_DW) - 1) : ((2 - NAlerts) * (2 - CLASS_DW)) + (((CLASS_DW - 1) + ((NAlerts - 1) * (2 - CLASS_DW))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))))))))))) + 1)] = reg2hw[811-:24];
	assign reg2hw_wrap[((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))))-:((((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))))) >= (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)))))) ? ((((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))))) - (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1))))))) + 1 : ((((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)))))) - (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))))))) + 1)] = {reg2hw[191] & (((reg2hw[186] | reg2hw[187]) | reg2hw[188]) | reg2hw[189]), reg2hw[383] & (((reg2hw[378] | reg2hw[379]) | reg2hw[380]) | reg2hw[381]), reg2hw[575] & (((reg2hw[570] | reg2hw[571]) | reg2hw[572]) | reg2hw[573]), reg2hw[767] & (((reg2hw[762] | reg2hw[763]) | reg2hw[764]) | reg2hw[765])};
	assign class_autolock_en = {reg2hw[190], reg2hw[382], reg2hw[574], reg2hw[766]};
	assign reg2hw_wrap[(((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)-:(((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)) >= ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)) - ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)) + 1 : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) - ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))) + 1)] = {reg2hw[186], reg2hw[187], reg2hw[188], reg2hw[189], reg2hw[378], reg2hw[379], reg2hw[380], reg2hw[381], reg2hw[570], reg2hw[571], reg2hw[572], reg2hw[573], reg2hw[762], reg2hw[763], reg2hw[764], reg2hw[765]};
	assign reg2hw_wrap[((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1-:((((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1) >= 0 ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) : 1 - (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))] = {reg2hw[179-:2], reg2hw[181-:2], reg2hw[183-:2], reg2hw[185-:2], reg2hw[371-:2], reg2hw[373-:2], reg2hw[375-:2], reg2hw[377-:2], reg2hw[563-:2], reg2hw[565-:2], reg2hw[567-:2], reg2hw[569-:2], reg2hw[755-:2], reg2hw[757-:2], reg2hw[759-:2], reg2hw[761-:2]};
	assign reg2hw_wrap[((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))))-:((((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))))) >= ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1))))) ? ((((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))))) - ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)))))) + 1 : (((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1))))) - (((N_CLASSES - 1) >= 0 ? N_CLASSES : 2 - N_CLASSES) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))))) + 1)] = {reg2hw[177] & reg2hw[176], reg2hw[369] & reg2hw[368], reg2hw[561] & reg2hw[560], reg2hw[753] & reg2hw[752]};
	assign reg2hw_wrap[(((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))-:(((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))) >= ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)))) ? (((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))) - ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1))))) + 1 : (((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)))) - ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))))) + 1)] = {reg2hw[175-:16], reg2hw[367-:16], reg2hw[559-:16], reg2hw[751-:16]};
	assign reg2hw_wrap[(((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))-:(((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))) >= (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1))) ? (((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))) - (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)))) + 1 : ((((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1))) - ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))))) + 1)] = {reg2hw[159-:32], reg2hw[351-:32], reg2hw[543-:32], reg2hw[735-:32]};
	assign reg2hw_wrap[((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))-:((((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))) >= ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)) ? ((((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1))) - ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1))) + 1 : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1)) - (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) : ((EscCntDw - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw : (EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw)))) - (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) ? ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) * (2 - EscCntDw))) - 1)) : ((EscCntDw - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * EscCntDw) + ((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * EscCntDw) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? 0 : N_PHASES - 1) : ((N_PHASES - 1) >= 0 ? (N_CLASSES - 1) * N_PHASES : (N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES)))) - ((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1)))) + 1) * (2 - EscCntDw)) + (((EscCntDw - 1) + (((N_CLASSES - 1) >= 0 ? ((N_PHASES - 1) >= 0 ? (N_CLASSES * N_PHASES) + -1 : (N_CLASSES * (2 - N_PHASES)) + ((N_PHASES - 1) - 1)) : ((N_PHASES - 1) >= 0 ? ((2 - N_CLASSES) * N_PHASES) + (((N_CLASSES - 1) * N_PHASES) - 1) : ((2 - N_CLASSES) * (2 - N_PHASES)) + (((N_PHASES - 1) + ((N_CLASSES - 1) * (2 - N_PHASES))) - 1))) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) + (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) >= (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) ? ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))))) + 1 : ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) : ((PHASE_DW - 1) >= 0 ? ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW : (PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW)))) - (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) ? ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) * (2 - PHASE_DW))) - 1)) : ((PHASE_DW - 1) >= 0 ? (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * PHASE_DW) + ((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * PHASE_DW) - 1) : (((((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? 0 : N_ESC_SEV - 1) : ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES - 1) * N_ESC_SEV : (N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV)))) - ((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1)))) + 1) * (2 - PHASE_DW)) + (((PHASE_DW - 1) + (((N_CLASSES - 1) >= 0 ? ((N_ESC_SEV - 1) >= 0 ? (N_CLASSES * N_ESC_SEV) + -1 : (N_CLASSES * (2 - N_ESC_SEV)) + ((N_ESC_SEV - 1) - 1)) : ((N_ESC_SEV - 1) >= 0 ? ((2 - N_CLASSES) * N_ESC_SEV) + (((N_CLASSES - 1) * N_ESC_SEV) - 1) : ((2 - N_CLASSES) * (2 - N_ESC_SEV)) + (((N_ESC_SEV - 1) + ((N_CLASSES - 1) * (2 - N_ESC_SEV))) - 1))) * (2 - PHASE_DW))) - 1)))) + 1) + -1)))) + 1)] = {reg2hw[31-:32], reg2hw[63-:32], reg2hw[95-:32], reg2hw[127-:32], reg2hw[223-:32], reg2hw[255-:32], reg2hw[287-:32], reg2hw[319-:32], reg2hw[415-:32], reg2hw[447-:32], reg2hw[479-:32], reg2hw[511-:32], reg2hw[607-:32], reg2hw[639-:32], reg2hw[671-:32], reg2hw[703-:32]};
	generate
		for (k = 0; k < NAlerts; k = k + 1) begin : gen_alert_cause_dump
			assign crashdump_o[((NAlerts - 1) >= 0 ? (((NAlerts - 1) >= 0 ? NAlerts : 2 - NAlerts) + (((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))))) - ((NAlerts - 1) - k) : (((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1)))) + (0 - k))] = reg2hw[784 + k];
		end
	endgenerate
	generate
		for (k = 0; k < N_LOC_ALERT; k = k + 1) begin : gen_loc_alert_cause_dump
			assign crashdump_o[((N_LOC_ALERT - 1) >= 0 ? (((N_LOC_ALERT - 1) >= 0 ? N_LOC_ALERT : 2 - N_LOC_ALERT) + ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1)))) - ((N_LOC_ALERT - 1) - k) : ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1))) + (0 - k))] = reg2hw[768 + k];
		end
	endgenerate
	assign crashdump_o[(((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))-:(((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))) >= ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1)) ? (((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))) - ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1))) + 1 : (((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1)) - ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1)))) + 1)] = hw2reg_wrap[(((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))-:(((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))) >= ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1)) ? (((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))) - ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1))) + 1 : (((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1)) - ((((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? 0 : AccuCntDw - 1) : ((AccuCntDw - 1) >= 0 ? (N_CLASSES - 1) * AccuCntDw : (AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((AccuCntDw - 1) >= 0 ? (N_CLASSES * AccuCntDw) + -1 : (N_CLASSES * (2 - AccuCntDw)) + ((AccuCntDw - 1) - 1)) : ((AccuCntDw - 1) >= 0 ? ((2 - N_CLASSES) * AccuCntDw) + (((N_CLASSES - 1) * AccuCntDw) - 1) : ((2 - N_CLASSES) * (2 - AccuCntDw)) + (((AccuCntDw - 1) + ((N_CLASSES - 1) * (2 - AccuCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1)))) + 1)];
	assign crashdump_o[(((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1)-:(((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1)) >= (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) ? (((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1)) - (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1)) + 1 : ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) - ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))) + 1)] = hw2reg_wrap[(((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1)-:(((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1)) >= (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) ? (((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1)) - (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1)) + 1 : ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) - ((((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) >= ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) ? (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))))) + 1 : (((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? 0 : EscCntDw - 1) : ((EscCntDw - 1) >= 0 ? (N_CLASSES - 1) * EscCntDw : (EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw)))) - ((N_CLASSES - 1) >= 0 ? ((EscCntDw - 1) >= 0 ? (N_CLASSES * EscCntDw) + -1 : (N_CLASSES * (2 - EscCntDw)) + ((EscCntDw - 1) - 1)) : ((EscCntDw - 1) >= 0 ? ((2 - N_CLASSES) * EscCntDw) + (((N_CLASSES - 1) * EscCntDw) - 1) : ((2 - N_CLASSES) * (2 - EscCntDw)) + (((EscCntDw - 1) + ((N_CLASSES - 1) * (2 - EscCntDw))) - 1)))) + 1) + ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))) + 1)];
	assign crashdump_o[(((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1-:(((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1) >= 0 ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) : 1 - ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))] = hw2reg_wrap[(((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1-:(((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1) >= 0 ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) : 1 - ((((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) >= ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) ? (((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1)) - ((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3)) + 1 : (((N_CLASSES - 1) >= 0 ? 0 : (N_CLASSES - 1) * 3) - ((N_CLASSES - 1) >= 0 ? (N_CLASSES * 3) + -1 : ((2 - N_CLASSES) * 3) + (((N_CLASSES - 1) * 3) - 1))) + 1) + -1))];
endmodule
