(* CLASS="output" *)
module VPR_OPAD(outpad);
    input  wire outpad;

endmodule
