(* whitebox *)
module CE_USED(CE, CE_OUT);
    input wire CE;
    output wire CE_OUT;

    assign CE_OUT = CE;
endmodule
