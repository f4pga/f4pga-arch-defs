(* blackbox *)
module LOGICBOX (I, O);
	input wire I;
	output wire O;
endmodule
