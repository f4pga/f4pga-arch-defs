module progmem
(
// Closk & reset
input  wire         clk,
input  wire         rstn,

// PicoRV32 bus interface
input  wire         valid,
output wire         ready,
input  wire [31:0]  addr,
output wire [31:0]  rdata
);

// ============================================================================

localparam  MEM_SIZE_BITS   = 10; // In 32-bit words
localparam  MEM_SIZE        = 1 << MEM_SIZE_BITS;
localparam  MEM_ADDR_MASK   = 32'h0010_0000;

// ============================================================================

wire [MEM_SIZE_BITS-1:0]    mem_addr;
reg  [31:0]                 mem_data;

always @(posedge clk)
    case (mem_addr)

    'h0000: mem_data <= 32'h00000093;
    'h0001: mem_data <= 32'h00000193;
    'h0002: mem_data <= 32'h00000213;
    'h0003: mem_data <= 32'h00000293;
    'h0004: mem_data <= 32'h00000313;
    'h0005: mem_data <= 32'h00000393;
    'h0006: mem_data <= 32'h00000413;
    'h0007: mem_data <= 32'h00000493;
    'h0008: mem_data <= 32'h00000513;
    'h0009: mem_data <= 32'h00000593;
    'h000A: mem_data <= 32'h00000613;
    'h000B: mem_data <= 32'h00000693;
    'h000C: mem_data <= 32'h00000713;
    'h000D: mem_data <= 32'h00000793;
    'h000E: mem_data <= 32'h00000813;
    'h000F: mem_data <= 32'h00000893;
    'h0010: mem_data <= 32'h00000913;
    'h0011: mem_data <= 32'h00000993;
    'h0012: mem_data <= 32'h00000A13;
    'h0013: mem_data <= 32'h00000A93;
    'h0014: mem_data <= 32'h00000B13;
    'h0015: mem_data <= 32'h00000B93;
    'h0016: mem_data <= 32'h00000C13;
    'h0017: mem_data <= 32'h00000C93;
    'h0018: mem_data <= 32'h00000D13;
    'h0019: mem_data <= 32'h00000D93;
    'h001A: mem_data <= 32'h00000E13;
    'h001B: mem_data <= 32'h00000E93;
    'h001C: mem_data <= 32'h00000F13;
    'h001D: mem_data <= 32'h00000F93;
    'h001E: mem_data <= 32'h03000537;
    'h001F: mem_data <= 32'h00100593;
    'h0020: mem_data <= 32'h00B52023;
    'h0021: mem_data <= 32'h00000513;
    'h0022: mem_data <= 32'h00A52023;
    'h0023: mem_data <= 32'h00450513;
    'h0024: mem_data <= 32'hFE254CE3;
    'h0025: mem_data <= 32'h03000537;
    'h0026: mem_data <= 32'h00300593;
    'h0027: mem_data <= 32'h00B52023;
    'h0028: mem_data <= 32'h00001517;
    'h0029: mem_data <= 32'hB4050513;
    'h002A: mem_data <= 32'h00000593;
    'h002B: mem_data <= 32'h00000613;
    'h002C: mem_data <= 32'h00C5DC63;
    'h002D: mem_data <= 32'h00052683;
    'h002E: mem_data <= 32'h00D5A023;
    'h002F: mem_data <= 32'h00450513;
    'h0030: mem_data <= 32'h00458593;
    'h0031: mem_data <= 32'hFEC5C8E3;
    'h0032: mem_data <= 32'h03000537;
    'h0033: mem_data <= 32'h00700593;
    'h0034: mem_data <= 32'h00B52023;
    'h0035: mem_data <= 32'h00000513;
    'h0036: mem_data <= 32'h00000593;
    'h0037: mem_data <= 32'h00B55863;
    'h0038: mem_data <= 32'h00052023;
    'h0039: mem_data <= 32'h00450513;
    'h003A: mem_data <= 32'hFEB54CE3;
    'h003B: mem_data <= 32'h03000537;
    'h003C: mem_data <= 32'h00F00593;
    'h003D: mem_data <= 32'h00B52023;
    'h003E: mem_data <= 32'h015000EF;
    'h003F: mem_data <= 32'h0000006F;
    'h0040: mem_data <= 32'h020002B7;
    'h0041: mem_data <= 32'h12000313;
    'h0042: mem_data <= 32'h00629023;
    'h0043: mem_data <= 32'h000281A3;
    'h0044: mem_data <= 32'h02060863;
    'h0045: mem_data <= 32'h00800F13;
    'h0046: mem_data <= 32'h0FF67393;
    'h0047: mem_data <= 32'h0073DE93;
    'h0048: mem_data <= 32'h01D28023;
    'h0049: mem_data <= 32'h010EEE93;
    'h004A: mem_data <= 32'h01D28023;
    'h004B: mem_data <= 32'h00139393;
    'h004C: mem_data <= 32'h0FF3F393;
    'h004D: mem_data <= 32'hFFFF0F13;
    'h004E: mem_data <= 32'hFE0F12E3;
    'h004F: mem_data <= 32'h00628023;
    'h0050: mem_data <= 32'h04058663;
    'h0051: mem_data <= 32'h00800F13;
    'h0052: mem_data <= 32'h00054383;
    'h0053: mem_data <= 32'h0073DE93;
    'h0054: mem_data <= 32'h01D28023;
    'h0055: mem_data <= 32'h010EEE93;
    'h0056: mem_data <= 32'h01D28023;
    'h0057: mem_data <= 32'h0002CE83;
    'h0058: mem_data <= 32'h002EFE93;
    'h0059: mem_data <= 32'h001EDE93;
    'h005A: mem_data <= 32'h00139393;
    'h005B: mem_data <= 32'h01D3E3B3;
    'h005C: mem_data <= 32'h0FF3F393;
    'h005D: mem_data <= 32'hFFFF0F13;
    'h005E: mem_data <= 32'hFC0F1AE3;
    'h005F: mem_data <= 32'h00750023;
    'h0060: mem_data <= 32'h00150513;
    'h0061: mem_data <= 32'hFFF58593;
    'h0062: mem_data <= 32'hFB9FF06F;
    'h0063: mem_data <= 32'h08000313;
    'h0064: mem_data <= 32'h006281A3;
    'h0065: mem_data <= 32'h00008067;
    'h0066: mem_data <= 32'hFE010113;
    'h0067: mem_data <= 32'h00112E23;
    'h0068: mem_data <= 32'h00812C23;
    'h0069: mem_data <= 32'h02010413;
    'h006A: mem_data <= 32'h00050793;
    'h006B: mem_data <= 32'hFEF407A3;
    'h006C: mem_data <= 32'hFEF44703;
    'h006D: mem_data <= 32'h00A00793;
    'h006E: mem_data <= 32'h00F71663;
    'h006F: mem_data <= 32'h00D00513;
    'h0070: mem_data <= 32'hFD9FF0EF;
    'h0071: mem_data <= 32'h020007B7;
    'h0072: mem_data <= 32'h00878793;
    'h0073: mem_data <= 32'hFEF44703;
    'h0074: mem_data <= 32'h00E7A023;
    'h0075: mem_data <= 32'h00000013;
    'h0076: mem_data <= 32'h01C12083;
    'h0077: mem_data <= 32'h01812403;
    'h0078: mem_data <= 32'h02010113;
    'h0079: mem_data <= 32'h00008067;
    'h007A: mem_data <= 32'hFE010113;
    'h007B: mem_data <= 32'h00112E23;
    'h007C: mem_data <= 32'h00812C23;
    'h007D: mem_data <= 32'h02010413;
    'h007E: mem_data <= 32'hFEA42623;
    'h007F: mem_data <= 32'h01C0006F;
    'h0080: mem_data <= 32'hFEC42783;
    'h0081: mem_data <= 32'h00178713;
    'h0082: mem_data <= 32'hFEE42623;
    'h0083: mem_data <= 32'h0007C783;
    'h0084: mem_data <= 32'h00078513;
    'h0085: mem_data <= 32'hF85FF0EF;
    'h0086: mem_data <= 32'hFEC42783;
    'h0087: mem_data <= 32'h0007C783;
    'h0088: mem_data <= 32'hFE0790E3;
    'h0089: mem_data <= 32'h00000013;
    'h008A: mem_data <= 32'h01C12083;
    'h008B: mem_data <= 32'h01812403;
    'h008C: mem_data <= 32'h02010113;
    'h008D: mem_data <= 32'h00008067;
    'h008E: mem_data <= 32'hFD010113;
    'h008F: mem_data <= 32'h02112623;
    'h0090: mem_data <= 32'h02812423;
    'h0091: mem_data <= 32'h03010413;
    'h0092: mem_data <= 32'hFCA42E23;
    'h0093: mem_data <= 32'hFCB42C23;
    'h0094: mem_data <= 32'h00700793;
    'h0095: mem_data <= 32'hFEF42623;
    'h0096: mem_data <= 32'h06C0006F;
    'h0097: mem_data <= 32'hFEC42783;
    'h0098: mem_data <= 32'h00279793;
    'h0099: mem_data <= 32'hFDC42703;
    'h009A: mem_data <= 32'h00F757B3;
    'h009B: mem_data <= 32'h00F7F713;
    'h009C: mem_data <= 32'h001017B7;
    'h009D: mem_data <= 32'hA8078793;
    'h009E: mem_data <= 32'h00F707B3;
    'h009F: mem_data <= 32'h0007C783;
    'h00A0: mem_data <= 32'hFEF405A3;
    'h00A1: mem_data <= 32'hFEB44703;
    'h00A2: mem_data <= 32'h03000793;
    'h00A3: mem_data <= 32'h00F71863;
    'h00A4: mem_data <= 32'hFEC42703;
    'h00A5: mem_data <= 32'hFD842783;
    'h00A6: mem_data <= 32'h00F75E63;
    'h00A7: mem_data <= 32'hFEB44783;
    'h00A8: mem_data <= 32'h00078513;
    'h00A9: mem_data <= 32'hEF5FF0EF;
    'h00AA: mem_data <= 32'hFEC42783;
    'h00AB: mem_data <= 32'hFCF42C23;
    'h00AC: mem_data <= 32'h0080006F;
    'h00AD: mem_data <= 32'h00000013;
    'h00AE: mem_data <= 32'hFEC42783;
    'h00AF: mem_data <= 32'hFFF78793;
    'h00B0: mem_data <= 32'hFEF42623;
    'h00B1: mem_data <= 32'hFEC42783;
    'h00B2: mem_data <= 32'hF807DAE3;
    'h00B3: mem_data <= 32'h00000013;
    'h00B4: mem_data <= 32'h02C12083;
    'h00B5: mem_data <= 32'h02812403;
    'h00B6: mem_data <= 32'h03010113;
    'h00B7: mem_data <= 32'h00008067;
    'h00B8: mem_data <= 32'hFE010113;
    'h00B9: mem_data <= 32'h00112E23;
    'h00BA: mem_data <= 32'h00812C23;
    'h00BB: mem_data <= 32'h02010413;
    'h00BC: mem_data <= 32'hFEA42623;
    'h00BD: mem_data <= 32'hFEC42703;
    'h00BE: mem_data <= 32'h06300793;
    'h00BF: mem_data <= 32'h00E7FA63;
    'h00C0: mem_data <= 32'h001017B7;
    'h00C1: mem_data <= 32'hA9478513;
    'h00C2: mem_data <= 32'hEE1FF0EF;
    'h00C3: mem_data <= 32'h28C0006F;
    'h00C4: mem_data <= 32'hFEC42703;
    'h00C5: mem_data <= 32'h05900793;
    'h00C6: mem_data <= 32'h00E7FE63;
    'h00C7: mem_data <= 32'h03900513;
    'h00C8: mem_data <= 32'hE79FF0EF;
    'h00C9: mem_data <= 32'hFEC42783;
    'h00CA: mem_data <= 32'hFA678793;
    'h00CB: mem_data <= 32'hFEF42623;
    'h00CC: mem_data <= 32'h1200006F;
    'h00CD: mem_data <= 32'hFEC42703;
    'h00CE: mem_data <= 32'h04F00793;
    'h00CF: mem_data <= 32'h00E7FE63;
    'h00D0: mem_data <= 32'h03800513;
    'h00D1: mem_data <= 32'hE55FF0EF;
    'h00D2: mem_data <= 32'hFEC42783;
    'h00D3: mem_data <= 32'hFB078793;
    'h00D4: mem_data <= 32'hFEF42623;
    'h00D5: mem_data <= 32'h0FC0006F;
    'h00D6: mem_data <= 32'hFEC42703;
    'h00D7: mem_data <= 32'h04500793;
    'h00D8: mem_data <= 32'h00E7FE63;
    'h00D9: mem_data <= 32'h03700513;
    'h00DA: mem_data <= 32'hE31FF0EF;
    'h00DB: mem_data <= 32'hFEC42783;
    'h00DC: mem_data <= 32'hFBA78793;
    'h00DD: mem_data <= 32'hFEF42623;
    'h00DE: mem_data <= 32'h0D80006F;
    'h00DF: mem_data <= 32'hFEC42703;
    'h00E0: mem_data <= 32'h03B00793;
    'h00E1: mem_data <= 32'h00E7FE63;
    'h00E2: mem_data <= 32'h03600513;
    'h00E3: mem_data <= 32'hE0DFF0EF;
    'h00E4: mem_data <= 32'hFEC42783;
    'h00E5: mem_data <= 32'hFC478793;
    'h00E6: mem_data <= 32'hFEF42623;
    'h00E7: mem_data <= 32'h0B40006F;
    'h00E8: mem_data <= 32'hFEC42703;
    'h00E9: mem_data <= 32'h03100793;
    'h00EA: mem_data <= 32'h00E7FE63;
    'h00EB: mem_data <= 32'h03500513;
    'h00EC: mem_data <= 32'hDE9FF0EF;
    'h00ED: mem_data <= 32'hFEC42783;
    'h00EE: mem_data <= 32'hFCE78793;
    'h00EF: mem_data <= 32'hFEF42623;
    'h00F0: mem_data <= 32'h0900006F;
    'h00F1: mem_data <= 32'hFEC42703;
    'h00F2: mem_data <= 32'h02700793;
    'h00F3: mem_data <= 32'h00E7FE63;
    'h00F4: mem_data <= 32'h03400513;
    'h00F5: mem_data <= 32'hDC5FF0EF;
    'h00F6: mem_data <= 32'hFEC42783;
    'h00F7: mem_data <= 32'hFD878793;
    'h00F8: mem_data <= 32'hFEF42623;
    'h00F9: mem_data <= 32'h06C0006F;
    'h00FA: mem_data <= 32'hFEC42703;
    'h00FB: mem_data <= 32'h01D00793;
    'h00FC: mem_data <= 32'h00E7FE63;
    'h00FD: mem_data <= 32'h03300513;
    'h00FE: mem_data <= 32'hDA1FF0EF;
    'h00FF: mem_data <= 32'hFEC42783;
    'h0100: mem_data <= 32'hFE278793;
    'h0101: mem_data <= 32'hFEF42623;
    'h0102: mem_data <= 32'h0480006F;
    'h0103: mem_data <= 32'hFEC42703;
    'h0104: mem_data <= 32'h01300793;
    'h0105: mem_data <= 32'h00E7FE63;
    'h0106: mem_data <= 32'h03200513;
    'h0107: mem_data <= 32'hD7DFF0EF;
    'h0108: mem_data <= 32'hFEC42783;
    'h0109: mem_data <= 32'hFEC78793;
    'h010A: mem_data <= 32'hFEF42623;
    'h010B: mem_data <= 32'h0240006F;
    'h010C: mem_data <= 32'hFEC42703;
    'h010D: mem_data <= 32'h00900793;
    'h010E: mem_data <= 32'h00E7FC63;
    'h010F: mem_data <= 32'h03100513;
    'h0110: mem_data <= 32'hD59FF0EF;
    'h0111: mem_data <= 32'hFEC42783;
    'h0112: mem_data <= 32'hFF678793;
    'h0113: mem_data <= 32'hFEF42623;
    'h0114: mem_data <= 32'hFEC42703;
    'h0115: mem_data <= 32'h00800793;
    'h0116: mem_data <= 32'h00E7FE63;
    'h0117: mem_data <= 32'h03900513;
    'h0118: mem_data <= 32'hD39FF0EF;
    'h0119: mem_data <= 32'hFEC42783;
    'h011A: mem_data <= 32'hFF778793;
    'h011B: mem_data <= 32'hFEF42623;
    'h011C: mem_data <= 32'h1280006F;
    'h011D: mem_data <= 32'hFEC42703;
    'h011E: mem_data <= 32'h00700793;
    'h011F: mem_data <= 32'h00E7FE63;
    'h0120: mem_data <= 32'h03800513;
    'h0121: mem_data <= 32'hD15FF0EF;
    'h0122: mem_data <= 32'hFEC42783;
    'h0123: mem_data <= 32'hFF878793;
    'h0124: mem_data <= 32'hFEF42623;
    'h0125: mem_data <= 32'h1040006F;
    'h0126: mem_data <= 32'hFEC42703;
    'h0127: mem_data <= 32'h00600793;
    'h0128: mem_data <= 32'h00E7FE63;
    'h0129: mem_data <= 32'h03700513;
    'h012A: mem_data <= 32'hCF1FF0EF;
    'h012B: mem_data <= 32'hFEC42783;
    'h012C: mem_data <= 32'hFF978793;
    'h012D: mem_data <= 32'hFEF42623;
    'h012E: mem_data <= 32'h0E00006F;
    'h012F: mem_data <= 32'hFEC42703;
    'h0130: mem_data <= 32'h00500793;
    'h0131: mem_data <= 32'h00E7FE63;
    'h0132: mem_data <= 32'h03600513;
    'h0133: mem_data <= 32'hCCDFF0EF;
    'h0134: mem_data <= 32'hFEC42783;
    'h0135: mem_data <= 32'hFFA78793;
    'h0136: mem_data <= 32'hFEF42623;
    'h0137: mem_data <= 32'h0BC0006F;
    'h0138: mem_data <= 32'hFEC42703;
    'h0139: mem_data <= 32'h00400793;
    'h013A: mem_data <= 32'h00E7FE63;
    'h013B: mem_data <= 32'h03500513;
    'h013C: mem_data <= 32'hCA9FF0EF;
    'h013D: mem_data <= 32'hFEC42783;
    'h013E: mem_data <= 32'hFFB78793;
    'h013F: mem_data <= 32'hFEF42623;
    'h0140: mem_data <= 32'h0980006F;
    'h0141: mem_data <= 32'hFEC42703;
    'h0142: mem_data <= 32'h00300793;
    'h0143: mem_data <= 32'h00E7FE63;
    'h0144: mem_data <= 32'h03400513;
    'h0145: mem_data <= 32'hC85FF0EF;
    'h0146: mem_data <= 32'hFEC42783;
    'h0147: mem_data <= 32'hFFC78793;
    'h0148: mem_data <= 32'hFEF42623;
    'h0149: mem_data <= 32'h0740006F;
    'h014A: mem_data <= 32'hFEC42703;
    'h014B: mem_data <= 32'h00200793;
    'h014C: mem_data <= 32'h00E7FE63;
    'h014D: mem_data <= 32'h03300513;
    'h014E: mem_data <= 32'hC61FF0EF;
    'h014F: mem_data <= 32'hFEC42783;
    'h0150: mem_data <= 32'hFFD78793;
    'h0151: mem_data <= 32'hFEF42623;
    'h0152: mem_data <= 32'h0500006F;
    'h0153: mem_data <= 32'hFEC42703;
    'h0154: mem_data <= 32'h00100793;
    'h0155: mem_data <= 32'h00E7FE63;
    'h0156: mem_data <= 32'h03200513;
    'h0157: mem_data <= 32'hC3DFF0EF;
    'h0158: mem_data <= 32'hFEC42783;
    'h0159: mem_data <= 32'hFFE78793;
    'h015A: mem_data <= 32'hFEF42623;
    'h015B: mem_data <= 32'h02C0006F;
    'h015C: mem_data <= 32'hFEC42783;
    'h015D: mem_data <= 32'h00078E63;
    'h015E: mem_data <= 32'h03100513;
    'h015F: mem_data <= 32'hC1DFF0EF;
    'h0160: mem_data <= 32'hFEC42783;
    'h0161: mem_data <= 32'hFFF78793;
    'h0162: mem_data <= 32'hFEF42623;
    'h0163: mem_data <= 32'h00C0006F;
    'h0164: mem_data <= 32'h03000513;
    'h0165: mem_data <= 32'hC05FF0EF;
    'h0166: mem_data <= 32'h01C12083;
    'h0167: mem_data <= 32'h01812403;
    'h0168: mem_data <= 32'h02010113;
    'h0169: mem_data <= 32'h00008067;
    'h016A: mem_data <= 32'hFD010113;
    'h016B: mem_data <= 32'h02112623;
    'h016C: mem_data <= 32'h02812423;
    'h016D: mem_data <= 32'h03010413;
    'h016E: mem_data <= 32'hFCA42E23;
    'h016F: mem_data <= 32'hFFF00793;
    'h0170: mem_data <= 32'hFEF42623;
    'h0171: mem_data <= 32'hC00027F3;
    'h0172: mem_data <= 32'hFEF42423;
    'h0173: mem_data <= 32'h030007B7;
    'h0174: mem_data <= 32'hFFF00713;
    'h0175: mem_data <= 32'h00E7A023;
    'h0176: mem_data <= 32'hFDC42783;
    'h0177: mem_data <= 32'h08078A63;
    'h0178: mem_data <= 32'hFDC42503;
    'h0179: mem_data <= 32'hC05FF0EF;
    'h017A: mem_data <= 32'h0880006F;
    'h017B: mem_data <= 32'hC00027F3;
    'h017C: mem_data <= 32'hFEF42223;
    'h017D: mem_data <= 32'hFE442703;
    'h017E: mem_data <= 32'hFE842783;
    'h017F: mem_data <= 32'h40F707B3;
    'h0180: mem_data <= 32'hFEF42023;
    'h0181: mem_data <= 32'hFE042703;
    'h0182: mem_data <= 32'h00B727B7;
    'h0183: mem_data <= 32'hB0078793;
    'h0184: mem_data <= 32'h04E7F863;
    'h0185: mem_data <= 32'hFDC42783;
    'h0186: mem_data <= 32'h00078663;
    'h0187: mem_data <= 32'hFDC42503;
    'h0188: mem_data <= 32'hBC9FF0EF;
    'h0189: mem_data <= 32'hFE442783;
    'h018A: mem_data <= 32'hFEF42423;
    'h018B: mem_data <= 32'h030007B7;
    'h018C: mem_data <= 32'h0007A783;
    'h018D: mem_data <= 32'h00179713;
    'h018E: mem_data <= 32'h030007B7;
    'h018F: mem_data <= 32'h0007A783;
    'h0190: mem_data <= 32'h0017D793;
    'h0191: mem_data <= 32'h0017F793;
    'h0192: mem_data <= 32'h0017B793;
    'h0193: mem_data <= 32'h0FF7F793;
    'h0194: mem_data <= 32'h00078693;
    'h0195: mem_data <= 32'h030007B7;
    'h0196: mem_data <= 32'h00D76733;
    'h0197: mem_data <= 32'h00E7A023;
    'h0198: mem_data <= 32'h020007B7;
    'h0199: mem_data <= 32'h00878793;
    'h019A: mem_data <= 32'h0007A783;
    'h019B: mem_data <= 32'hFEF42623;
    'h019C: mem_data <= 32'hFEC42703;
    'h019D: mem_data <= 32'hFFF00793;
    'h019E: mem_data <= 32'hF6F70AE3;
    'h019F: mem_data <= 32'h030007B7;
    'h01A0: mem_data <= 32'h0007A023;
    'h01A1: mem_data <= 32'hFEC42783;
    'h01A2: mem_data <= 32'h0FF7F793;
    'h01A3: mem_data <= 32'h00078513;
    'h01A4: mem_data <= 32'h02C12083;
    'h01A5: mem_data <= 32'h02812403;
    'h01A6: mem_data <= 32'h03010113;
    'h01A7: mem_data <= 32'h00008067;
    'h01A8: mem_data <= 32'hFF010113;
    'h01A9: mem_data <= 32'h00112623;
    'h01AA: mem_data <= 32'h00812423;
    'h01AB: mem_data <= 32'h01010413;
    'h01AC: mem_data <= 32'h00000513;
    'h01AD: mem_data <= 32'hEF5FF0EF;
    'h01AE: mem_data <= 32'h00050793;
    'h01AF: mem_data <= 32'h00078513;
    'h01B0: mem_data <= 32'h00C12083;
    'h01B1: mem_data <= 32'h00812403;
    'h01B2: mem_data <= 32'h01010113;
    'h01B3: mem_data <= 32'h00008067;
    'h01B4: mem_data <= 32'hEB010113;
    'h01B5: mem_data <= 32'h14112623;
    'h01B6: mem_data <= 32'h14812423;
    'h01B7: mem_data <= 32'h15010413;
    'h01B8: mem_data <= 32'h00050793;
    'h01B9: mem_data <= 32'hEAB42C23;
    'h01BA: mem_data <= 32'hEAF40FA3;
    'h01BB: mem_data <= 32'hEC040793;
    'h01BC: mem_data <= 32'hFCF42A23;
    'h01BD: mem_data <= 32'h12B9B7B7;
    'h01BE: mem_data <= 32'h0A178793;
    'h01BF: mem_data <= 32'hFEF42623;
    'h01C0: mem_data <= 32'hC00027F3;
    'h01C1: mem_data <= 32'hFCF42823;
    'h01C2: mem_data <= 32'hC02027F3;
    'h01C3: mem_data <= 32'hFCF42623;
    'h01C4: mem_data <= 32'hFE042423;
    'h01C5: mem_data <= 32'h1200006F;
    'h01C6: mem_data <= 32'hFE042223;
    'h01C7: mem_data <= 32'h0640006F;
    'h01C8: mem_data <= 32'hFEC42783;
    'h01C9: mem_data <= 32'h00D79793;
    'h01CA: mem_data <= 32'hFEC42703;
    'h01CB: mem_data <= 32'h00F747B3;
    'h01CC: mem_data <= 32'hFEF42623;
    'h01CD: mem_data <= 32'hFEC42783;
    'h01CE: mem_data <= 32'h0117D793;
    'h01CF: mem_data <= 32'hFEC42703;
    'h01D0: mem_data <= 32'h00F747B3;
    'h01D1: mem_data <= 32'hFEF42623;
    'h01D2: mem_data <= 32'hFEC42783;
    'h01D3: mem_data <= 32'h00579793;
    'h01D4: mem_data <= 32'hFEC42703;
    'h01D5: mem_data <= 32'h00F747B3;
    'h01D6: mem_data <= 32'hFEF42623;
    'h01D7: mem_data <= 32'hFEC42783;
    'h01D8: mem_data <= 32'h0FF7F713;
    'h01D9: mem_data <= 32'hFE442783;
    'h01DA: mem_data <= 32'hFF040693;
    'h01DB: mem_data <= 32'h00F687B3;
    'h01DC: mem_data <= 32'hECE78823;
    'h01DD: mem_data <= 32'hFE442783;
    'h01DE: mem_data <= 32'h00178793;
    'h01DF: mem_data <= 32'hFEF42223;
    'h01E0: mem_data <= 32'hFE442703;
    'h01E1: mem_data <= 32'h0FF00793;
    'h01E2: mem_data <= 32'hF8E7DCE3;
    'h01E3: mem_data <= 32'hFE042023;
    'h01E4: mem_data <= 32'hFC042E23;
    'h01E5: mem_data <= 32'h0440006F;
    'h01E6: mem_data <= 32'hFE042783;
    'h01E7: mem_data <= 32'hFF040713;
    'h01E8: mem_data <= 32'h00F707B3;
    'h01E9: mem_data <= 32'hED07C783;
    'h01EA: mem_data <= 32'h02078263;
    'h01EB: mem_data <= 32'hFDC42783;
    'h01EC: mem_data <= 32'h00178713;
    'h01ED: mem_data <= 32'hFCE42E23;
    'h01EE: mem_data <= 32'hFE042703;
    'h01EF: mem_data <= 32'h0FF77713;
    'h01F0: mem_data <= 32'hFF040693;
    'h01F1: mem_data <= 32'h00F687B3;
    'h01F2: mem_data <= 32'hECE78823;
    'h01F3: mem_data <= 32'hFE042783;
    'h01F4: mem_data <= 32'h00178793;
    'h01F5: mem_data <= 32'hFEF42023;
    'h01F6: mem_data <= 32'hFE042703;
    'h01F7: mem_data <= 32'h0FF00793;
    'h01F8: mem_data <= 32'hFAE7DCE3;
    'h01F9: mem_data <= 32'hFC042C23;
    'h01FA: mem_data <= 32'hFC042023;
    'h01FB: mem_data <= 32'h0300006F;
    'h01FC: mem_data <= 32'hFD842783;
    'h01FD: mem_data <= 32'h00279793;
    'h01FE: mem_data <= 32'hFD442703;
    'h01FF: mem_data <= 32'h00F707B3;
    'h0200: mem_data <= 32'h0007A783;
    'h0201: mem_data <= 32'hFEC42703;
    'h0202: mem_data <= 32'h00F747B3;
    'h0203: mem_data <= 32'hFEF42623;
    'h0204: mem_data <= 32'hFD842783;
    'h0205: mem_data <= 32'h00178793;
    'h0206: mem_data <= 32'hFCF42C23;
    'h0207: mem_data <= 32'hFD842703;
    'h0208: mem_data <= 32'h03F00793;
    'h0209: mem_data <= 32'hFCE7D6E3;
    'h020A: mem_data <= 32'hFE842783;
    'h020B: mem_data <= 32'h00178793;
    'h020C: mem_data <= 32'hFEF42423;
    'h020D: mem_data <= 32'hFE842703;
    'h020E: mem_data <= 32'h01300793;
    'h020F: mem_data <= 32'hECE7DEE3;
    'h0210: mem_data <= 32'hC00027F3;
    'h0211: mem_data <= 32'hFCF42423;
    'h0212: mem_data <= 32'hC02027F3;
    'h0213: mem_data <= 32'hFCF42223;
    'h0214: mem_data <= 32'hEBF44783;
    'h0215: mem_data <= 32'h06078E63;
    'h0216: mem_data <= 32'h001017B7;
    'h0217: mem_data <= 32'hA9C78513;
    'h0218: mem_data <= 32'h989FF0EF;
    'h0219: mem_data <= 32'hFC842703;
    'h021A: mem_data <= 32'hFD042783;
    'h021B: mem_data <= 32'h40F707B3;
    'h021C: mem_data <= 32'h00800593;
    'h021D: mem_data <= 32'h00078513;
    'h021E: mem_data <= 32'h9C1FF0EF;
    'h021F: mem_data <= 32'h00A00513;
    'h0220: mem_data <= 32'h919FF0EF;
    'h0221: mem_data <= 32'h001017B7;
    'h0222: mem_data <= 32'hAA878513;
    'h0223: mem_data <= 32'h95DFF0EF;
    'h0224: mem_data <= 32'hFC442703;
    'h0225: mem_data <= 32'hFCC42783;
    'h0226: mem_data <= 32'h40F707B3;
    'h0227: mem_data <= 32'h00800593;
    'h0228: mem_data <= 32'h00078513;
    'h0229: mem_data <= 32'h995FF0EF;
    'h022A: mem_data <= 32'h00A00513;
    'h022B: mem_data <= 32'h8EDFF0EF;
    'h022C: mem_data <= 32'h001017B7;
    'h022D: mem_data <= 32'hAB478513;
    'h022E: mem_data <= 32'h931FF0EF;
    'h022F: mem_data <= 32'h00800593;
    'h0230: mem_data <= 32'hFEC42503;
    'h0231: mem_data <= 32'h975FF0EF;
    'h0232: mem_data <= 32'h00A00513;
    'h0233: mem_data <= 32'h8CDFF0EF;
    'h0234: mem_data <= 32'hEB842783;
    'h0235: mem_data <= 32'h00078C63;
    'h0236: mem_data <= 32'hFC442703;
    'h0237: mem_data <= 32'hFCC42783;
    'h0238: mem_data <= 32'h40F70733;
    'h0239: mem_data <= 32'hEB842783;
    'h023A: mem_data <= 32'h00E7A023;
    'h023B: mem_data <= 32'hFC842703;
    'h023C: mem_data <= 32'hFD042783;
    'h023D: mem_data <= 32'h40F707B3;
    'h023E: mem_data <= 32'h00078513;
    'h023F: mem_data <= 32'h14C12083;
    'h0240: mem_data <= 32'h14812403;
    'h0241: mem_data <= 32'h15010113;
    'h0242: mem_data <= 32'h00008067;
    'h0243: mem_data <= 32'hFE010113;
    'h0244: mem_data <= 32'h00112E23;
    'h0245: mem_data <= 32'h00812C23;
    'h0246: mem_data <= 32'h02010413;
    'h0247: mem_data <= 32'h030007B7;
    'h0248: mem_data <= 32'h01F00713;
    'h0249: mem_data <= 32'h00E7A023;
    'h024A: mem_data <= 32'h020007B7;
    'h024B: mem_data <= 32'h00478793;
    'h024C: mem_data <= 32'h36400713;
    'h024D: mem_data <= 32'h00E7A023;
    'h024E: mem_data <= 32'h001017B7;
    'h024F: mem_data <= 32'hAC078513;
    'h0250: mem_data <= 32'h8A9FF0EF;
    'h0251: mem_data <= 32'h030007B7;
    'h0252: mem_data <= 32'h03F00713;
    'h0253: mem_data <= 32'h00E7A023;
    'h0254: mem_data <= 32'h030007B7;
    'h0255: mem_data <= 32'h07F00713;
    'h0256: mem_data <= 32'h00E7A023;
    'h0257: mem_data <= 32'h00000013;
    'h0258: mem_data <= 32'h001017B7;
    'h0259: mem_data <= 32'hACC78513;
    'h025A: mem_data <= 32'hC41FF0EF;
    'h025B: mem_data <= 32'h00050793;
    'h025C: mem_data <= 32'h00078713;
    'h025D: mem_data <= 32'h00D00793;
    'h025E: mem_data <= 32'hFEF714E3;
    'h025F: mem_data <= 32'h001017B7;
    'h0260: mem_data <= 32'hAE878513;
    'h0261: mem_data <= 32'h865FF0EF;
    'h0262: mem_data <= 32'h001017B7;
    'h0263: mem_data <= 32'hAEC78513;
    'h0264: mem_data <= 32'h859FF0EF;
    'h0265: mem_data <= 32'h001017B7;
    'h0266: mem_data <= 32'hB1478513;
    'h0267: mem_data <= 32'h84DFF0EF;
    'h0268: mem_data <= 32'h001017B7;
    'h0269: mem_data <= 32'hB3C78513;
    'h026A: mem_data <= 32'h841FF0EF;
    'h026B: mem_data <= 32'h001017B7;
    'h026C: mem_data <= 32'hB6078513;
    'h026D: mem_data <= 32'h835FF0EF;
    'h026E: mem_data <= 32'h001017B7;
    'h026F: mem_data <= 32'hB8878513;
    'h0270: mem_data <= 32'h829FF0EF;
    'h0271: mem_data <= 32'h001017B7;
    'h0272: mem_data <= 32'hAE878513;
    'h0273: mem_data <= 32'h81DFF0EF;
    'h0274: mem_data <= 32'h001017B7;
    'h0275: mem_data <= 32'hAE878513;
    'h0276: mem_data <= 32'h811FF0EF;
    'h0277: mem_data <= 32'h001017B7;
    'h0278: mem_data <= 32'hBB078513;
    'h0279: mem_data <= 32'h805FF0EF;
    'h027A: mem_data <= 32'h001017B7;
    'h027B: mem_data <= 32'hAE878513;
    'h027C: mem_data <= 32'hFF8FF0EF;
    'h027D: mem_data <= 32'h00A00793;
    'h027E: mem_data <= 32'hFEF42623;
    'h027F: mem_data <= 32'h0780006F;
    'h0280: mem_data <= 32'h001017B7;
    'h0281: mem_data <= 32'hBD478513;
    'h0282: mem_data <= 32'hFE0FF0EF;
    'h0283: mem_data <= 32'hC95FF0EF;
    'h0284: mem_data <= 32'h00050793;
    'h0285: mem_data <= 32'hFEF405A3;
    'h0286: mem_data <= 32'hFEB44703;
    'h0287: mem_data <= 32'h02000793;
    'h0288: mem_data <= 32'h00E7FE63;
    'h0289: mem_data <= 32'hFEB44703;
    'h028A: mem_data <= 32'h07E00793;
    'h028B: mem_data <= 32'h00E7E863;
    'h028C: mem_data <= 32'hFEB44783;
    'h028D: mem_data <= 32'h00078513;
    'h028E: mem_data <= 32'hF60FF0EF;
    'h028F: mem_data <= 32'h001017B7;
    'h0290: mem_data <= 32'hAE878513;
    'h0291: mem_data <= 32'hFA4FF0EF;
    'h0292: mem_data <= 32'hFEB44703;
    'h0293: mem_data <= 32'h03900793;
    'h0294: mem_data <= 32'h00F71C63;
    'h0295: mem_data <= 32'h00000593;
    'h0296: mem_data <= 32'h00100513;
    'h0297: mem_data <= 32'hC75FF0EF;
    'h0298: mem_data <= 32'h00000013;
    'h0299: mem_data <= 32'h0180006F;
    'h029A: mem_data <= 32'hFEC42783;
    'h029B: mem_data <= 32'hFFF78793;
    'h029C: mem_data <= 32'hFEF42623;
    'h029D: mem_data <= 32'hFEC42783;
    'h029E: mem_data <= 32'hF8F044E3;
    'h029F: mem_data <= 32'hF49FF06F;
    'h02A0: mem_data <= 32'h33323130;
    'h02A1: mem_data <= 32'h37363534;
    'h02A2: mem_data <= 32'h62613938;
    'h02A3: mem_data <= 32'h66656463;
    'h02A4: mem_data <= 32'h00000000;
    'h02A5: mem_data <= 32'h30313D3E;
    'h02A6: mem_data <= 32'h00000030;
    'h02A7: mem_data <= 32'h6C637943;
    'h02A8: mem_data <= 32'h203A7365;
    'h02A9: mem_data <= 32'h00007830;
    'h02AA: mem_data <= 32'h74736E49;
    'h02AB: mem_data <= 32'h203A736E;
    'h02AC: mem_data <= 32'h00007830;
    'h02AD: mem_data <= 32'h736B6843;
    'h02AE: mem_data <= 32'h203A6D75;
    'h02AF: mem_data <= 32'h00007830;
    'h02B0: mem_data <= 32'h746F6F42;
    'h02B1: mem_data <= 32'h2E676E69;
    'h02B2: mem_data <= 32'h00000A2E;
    'h02B3: mem_data <= 32'h73657250;
    'h02B4: mem_data <= 32'h4E452073;
    'h02B5: mem_data <= 32'h20524554;
    'h02B6: mem_data <= 32'h63206F74;
    'h02B7: mem_data <= 32'h69746E6F;
    'h02B8: mem_data <= 32'h2E65756E;
    'h02B9: mem_data <= 32'h00000A2E;
    'h02BA: mem_data <= 32'h0000000A;
    'h02BB: mem_data <= 32'h5F5F2020;
    'h02BC: mem_data <= 32'h20205F5F;
    'h02BD: mem_data <= 32'h2020205F;
    'h02BE: mem_data <= 32'h20202020;
    'h02BF: mem_data <= 32'h5F202020;
    'h02C0: mem_data <= 32'h205F5F5F;
    'h02C1: mem_data <= 32'h20202020;
    'h02C2: mem_data <= 32'h20202020;
    'h02C3: mem_data <= 32'h5F5F5F5F;
    'h02C4: mem_data <= 32'h0000000A;
    'h02C5: mem_data <= 32'h20207C20;
    'h02C6: mem_data <= 32'h285C205F;
    'h02C7: mem_data <= 32'h5F20295F;
    'h02C8: mem_data <= 32'h5F205F5F;
    'h02C9: mem_data <= 32'h202F5F5F;
    'h02CA: mem_data <= 32'h7C5F5F5F;
    'h02CB: mem_data <= 32'h5F5F2020;
    'h02CC: mem_data <= 32'h2F20205F;
    'h02CD: mem_data <= 32'h5F5F5F20;
    'h02CE: mem_data <= 32'h00000A7C;
    'h02CF: mem_data <= 32'h7C207C20;
    'h02D0: mem_data <= 32'h7C20295F;
    'h02D1: mem_data <= 32'h202F7C20;
    'h02D2: mem_data <= 32'h202F5F5F;
    'h02D3: mem_data <= 32'h5F5C205F;
    'h02D4: mem_data <= 32'h5C205F5F;
    'h02D5: mem_data <= 32'h5F202F20;
    'h02D6: mem_data <= 32'h207C5C20;
    'h02D7: mem_data <= 32'h00000A7C;
    'h02D8: mem_data <= 32'h20207C20;
    'h02D9: mem_data <= 32'h7C2F5F5F;
    'h02DA: mem_data <= 32'h28207C20;
    'h02DB: mem_data <= 32'h28207C5F;
    'h02DC: mem_data <= 32'h7C20295F;
    'h02DD: mem_data <= 32'h20295F5F;
    'h02DE: mem_data <= 32'h5F28207C;
    'h02DF: mem_data <= 32'h207C2029;
    'h02E0: mem_data <= 32'h5F5F5F7C;
    'h02E1: mem_data <= 32'h0000000A;
    'h02E2: mem_data <= 32'h7C5F7C20;
    'h02E3: mem_data <= 32'h7C202020;
    'h02E4: mem_data <= 32'h5F5C7C5F;
    'h02E5: mem_data <= 32'h5F5C5F5F;
    'h02E6: mem_data <= 32'h5F2F5F5F;
    'h02E7: mem_data <= 32'h2F5F5F5F;
    'h02E8: mem_data <= 32'h5F5F5C20;
    'h02E9: mem_data <= 32'h5C202F5F;
    'h02EA: mem_data <= 32'h5F5F5F5F;
    'h02EB: mem_data <= 32'h00000A7C;
    'h02EC: mem_data <= 32'h5B202020;
    'h02ED: mem_data <= 32'h52205D39;
    'h02EE: mem_data <= 32'h73206E75;
    'h02EF: mem_data <= 32'h6C706D69;
    'h02F0: mem_data <= 32'h69747369;
    'h02F1: mem_data <= 32'h65622063;
    'h02F2: mem_data <= 32'h6D68636E;
    'h02F3: mem_data <= 32'h0A6B7261;
    'h02F4: mem_data <= 32'h00000000;
    'h02F5: mem_data <= 32'h6D6D6F43;
    'h02F6: mem_data <= 32'h3E646E61;
    'h02F7: mem_data <= 32'h00000020;

    default:    mem_data <= 32'hDEADBEEF;

    endcase

// ============================================================================

reg o_ready;

always @(posedge clk or negedge rstn)
    if (!rstn)  o_ready <= 1'd0;
    else        o_ready <= valid && ((addr & MEM_ADDR_MASK) != 0);

// Output connectins
assign ready    = o_ready;
assign rdata    = mem_data;
assign mem_addr = addr[MEM_SIZE_BITS+1:2];

endmodule

