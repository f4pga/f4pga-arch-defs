(* whitebox *)
module SR_GND(SR_OUT);
    output wire SR_OUT;

    assign SR_OUT = 1;
endmodule
