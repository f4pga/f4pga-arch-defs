`define SEED 32'h94e264fd
