module top (
	input  clk,
	input [15:0] in,
	output [3:0] out
);
    DPRAM64D #(
        .INIT(64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010)
    ) ram3(
        .CLK(clk),
        .A(in[5:0]),
        .O6(out[3]),
        .DI1(in[14]),
        .WE(in[15])
    );
    DPRAM64C #(
        .INIT(64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010)
    ) ram4(
        .CLK(clk),
        .A(in[5:0]),
        .O6(out[2]),
        .DI1(in[13]),
        .WE(in[15])
    );

    DPRAM64B #(
        .INIT(64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010)
    ) ram1(
        .CLK(clk),
        .A(in[5:0]),
        .O6(out[1]),
        .DI1(in[12]),
        .WE(in[15])
    );
    DPRAM64A #(
        .INIT(64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010)
    ) ram2(
        .CLK(clk),
        .A(in[5:0]),
        .O6(out[0]),
        .DI1(in[11]),
        .WE(in[15])
    );
endmodule
